-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����X��V������6�8�!�%�+���Y����\��}��U���0�8�;�x�w�/����Ӷ��Y��N��<���c�`�_�x��)�M��Y����Q��^����x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��Yۅ�V��-�����=�u�4�<�9�1�>�������G��X�����:�_�x��;�����Y����A��=C�;���:�4�u�;�#�(����Y����A��'�����!�:�_�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���9K�g�����u��6�4�2�;�����Ƹ�VF��V�����u�0�<�4�8�s�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�=d�����,���y� �/�L�������v#��D�����6�d�c�{�;�f�Wϫ�ӯ��vH��Z�����1�4�9�_�w�.�W���ݶ��u��C*��6���3�6�0�!�y�1�L�������VF��P(�����;�9�0�<�6�2�W���s���3��V�����&��6�0�2�)����
����G6��D��ʓ�4�!�0��8�����������=N��Xʼ�u��8�=�$���������@l�T�����u��8�=�$�����Y����T��S��F���x�u�g�{�e�}��������X(��t��%���0�<�&�o�>�)����C����F�=�[��_�u�x�>�"�����
����]�������u�4�<�u�#�n����
����WF��Z��U���=�;�0�{�w�p�W���������DN�����"� �1�'�&�4�ϼ�
�Ư�V ��T�����0�<�!�<�"�4��ԜY����eF��p/�����6�4�2�&�6�9����	������T��U���!�<�u�4�3�>�������K��X�����!�'�0��8�8����,����l�T�����u��8�'�4�.��������	F��C����u�n�_�u�z�	��������\��E�����=�u�'�4�w�4�Ϫ�Ӕ��[��B��ʺ�u�:�3�u�%�<�}���TӀ����_N�����&�;�u�;�#�W�W�������!��t�����8�'�4�}��8����0����]�������|�'�!�'�w��:������U��C��U����!�:�3��<�6��� ۍ��V ��R�����6�o�<�!�0�/�W�������a'��1����1��6�4�2���������R
��T�����_��6�4�2�?��������P��Y�����4�:�u�&�]�}��������V��R�����'�4�}��2�;����
����V\��Y�����'�!�'�u���A������F��E�����0� �;�'�6�}�W���4�Г�\������h�u�:�=�%�}�I���^����F��P��U���<�}��0�1�8�>�������F�����ߊu�u�u�0�"�3����Y����p	��Q#�����n�u�u�0�$�;��������z��V ��U���|�!�0�_�w�}�W�������A��S��6���3�0�:�,�l�}�Wϻ�
���F�e�����'�,�o�u��8��������9F���U���_�u�u�0�"�3�%�������R��N��ʒ�!�:�3��6�����s����F��^��2���9��0�3�%�0����Q����U ��Z'�����0�u�;�0�2�t�����Ǝ�r+��h�����u�#�'�4�;�}��������JF��u<��F܊�u�h�}�!�2�.�J�������@F�I�\��u�7�2�;�w�}����:����~��Y�����h�e�u�=�9�W�W���Y����A��E��O����0�3�0�8�$���s���V
��QF������8�;�!�9�8�J��Y����9F�N�����;�'�4�u�j�6����4����J'��UךU���9�0�u�u�w�����8����\�\-�����8�'��!�l�}�Wϻ�ӏ��9F��� ����!�'��%�$�}����Ƌ�G'��t�����8�'�4�n�2�9�'�������\��g�����<�;�9�0�>�<���