-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����u
��������!�:�o��<�ϝ�����K��E������:�0�!�w�4����s����R��Y�����u�e�e�x�]�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���l�F��U��e��%�'�0�)�9�������z��E������'�:�4�>�3�Z����ƞ�T��<�����1�x�u�4�>�3�ϗ�
����V��'�����9��3�'�6�4���T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�CחX���u� �%�&�m�p�W���-����P��C��ʳ�<�x�9�%�"�4�Ϫ�Ӿ��Z��C��1���u�:�!�,�#�}��������G��T��ʰ�4�9�u�;�]�p����Ӗ��GK��Y�����;�8�u�=�#�4�W�������\F��Y
�X�߇x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�}��������RUךU���u�0�0�&�3�1����H����R
��=d�����,�"�'�n�w�(�ϩ��Ȝ�T(��C�����{�9�n�_�>�/����7����l�B�� ����{�6�8�8�8������ƓV��C��3���u�&�u�2�9�/����+����e��N�����2�6�o�u�g�t�}������9F������u��u�o�>�}������ƹF��[����u�u�;�&�3�1����s���P7�T�� ���!�
�:�<�w�`��������9F�d�����<� �0�1�%�>�(��������[��N���4�!�<� �2�9����&����_��QN����&�2�4�u�$�)�������u
��d�����!�6� �0�%�1����?����ZǑN����>�&�2�!�%�W�W�������p
����*���<�n�u�&�0�<�W����ƿ�W9��P�����x�=�:�
�>�8��ԜY����G�������}�0�0��;�g��������F��C��U���u�&�u�7�0�3�W����ƞ�@��V��E���=�;�'�!�%�}�G������A��E ��D��0�1�<�n�w�8�ϸ�����]F��R���ߠ7�2�;�_�w�p�#���Y����]F��S�����&��6�;�6�<��������R����ǳ�:�u�;�u�8�W�W���ƪ�\
�������1�9�4�1�;�$����Y����A��YN��ʅ��4�1���.����
���t��d��8���9�u�3�3�;�8��������F�G�����}��&�!�w�1�^���Yӄ��ZǻN��U���4�0�0�u�?�3�W���Y����bF�I�N���u�u�0�&�1�/����&����%��N���ߊu�u�u�u�1�>�Ϫ��Ư�Z�T*����<�n�u�u�w�8�Ϸ�B����������n�u�0�1�0�3����Y����`��z���ߠu�x�#�6�9�+������ƓF�9�����u�u�:�4�9�2�W���Ӈ����EN�����!�0�r�0�9�)����Y����[��X
��U���#�_�u�x�6�9����Y����_F����U���,�!�<�2��>�ϲ�����GHǻC�����
�:�4�;�6�/�}���T����X9��@��U���'�u�4�'�w�`�P�������R4��R������&�!�4�j�l�W�������l�V-��U��r�r�"�0�w���������a��C8��H��u�9�0�r�p�W�W������l��s-�����x�=�:�
�w��#ϵ�������D�����u�x�#�:�<�<�'�������F�A�������4�9�]�}�Z�������pF��\d��Xǣ�:�>�4��w�2�$�������P#��=N��X���:�
�u�u��}�Z¨�����7��fd��3����o����}�WϹ�������FךU���u���h�w�����Q����V��[G��U���<�u�7�!�m�}�G�ԜY�Ƽ�A��V�����u�u��u�i�<���Y���F�N��X���;�u�!�
�8�4�}���Y�Ə�aF������u�u�u�u�w�}�Z����ƿ�W9��P��U���u��u�h�w�1�[���Y���F�N��Xʼ�u�&�1�9�0�>�W���Yӥ��[�c�����2�6�6�;�{�}�ZϷ�Yӕ��l
��^ךU���u�u�u�k�4�q�W���Y���F�N�U���u�!�
�:�>�W�W���Y���X��fG�U���u�u�u�u�w�p�W���Y����_	��TdךU���0��'�u�1�6����/���A��R �����u�x�_�u�z�}�Z�������u"��(�����x�u�x�#�8�6�ϗ�0�ƣ�VǻC�U���=�:�
�u��}��������PN��R��\���x�u�x�#�8�6�ϝ�:��ƹK�C�����
�u����)�;���ۅ��l�C��Xǣ�:�>�4��4�W�W��Y�˺�\	��VN���ߊu�x�u��/�}�3���Y���F��R �����4�u�_�u�z�}�W���7���F��R ��U���<�u�7�!�m�}�G�ԜY���F��E�����_�u�x�u�w�}�;���GӲ��`��X	��]���&�!�y�u�z�4�Wϭ�����ZǻC�U���u�u�u�k��6�W���Y���F�N��U���<�u�&�1�;�:����T���F��rN��Kʁ�
�!��2�4�>���Y���F��N�����2�6�u�x�w�}�WϚ�Y���P"�N��U���u�u�u�u�w�p�W���Y����_	��Td��X���u�u��u�j�}�&��Y���F�N��U���x�u� �u�#�����s���9F���U���0�4�0��9�1�L���T���K��Y=��Oʼ�u��&�!�6�`�F�������GǻC�U���u�x�#�:�<�4�1���Y����9F�N��X���:�
�u���2��ԜY���K��X��ʅ���
�!��:�ǿ�����9F�N��X���:�
�u�u�;�W�W��Y�˺�\	��VN��U����1�:�<���^���T�����X��U����u�x�u�z�+����ӷ��bl�C��3���o���_�w�p�W�������PF��GN��U���u�u�u���}�Iϱ����K��YN�����h�r�r�u�z�}�WϮ��ơ�CF�N�U���u���h�w�2�$�������R4��R��U���u�;�u�!��2��ԜY���F�tN��H���9�y�u�u�w�}�W���Y���K��YN�����:�<�_�u�z�}�W���<���2��d�����}��|�u�w�}�ZϷ�Yӕ��l
��^ךU���u�u�u�u�w�c���Y���F�N��U���u�x�<�u�$�9�������F�N��U���k�6�|�u�w�}�W���Y���F�N��ʦ�1�9�2�6�w�p�}���T����T��E��U����!�_�u�z�}�Z¨�����@��h�����u�!�n�_�z�	�ϸ�����]��X�����&�4�6�0�<�(�W����ƹ�V��XN�����<�0�"�0�?�/����s����Z
��_�����u�:�<�<�3�}�'���
�ƨ�]A��C�����0�u�'� �3�4�Y���ԕ��[��=C����4�'�4�:�y�p�!�������S��Z�