-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����A��s�����;�!�#�1�z�}�����Ɔ�[��Z�����x�u�'�2�9�1�'�������c>��h[�@�߇x��!�o�e�}����K����KǶC�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�_�x��t�E��Y����A��CN�����4�u�;�!�"�8��������R��Yd�U���u�<�=�&��.����s����R��Y��<���'�8�;�&��)����Y����A��^��X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�}��)����@��:��ʳ�9�u�'�4�2�}��������@����ʳ�'�!�0�3�6�)����Y����^��E@חX���u�u�u�u��8��������TF��^��ʶ�8�:�0�u�1�<��������]�������<�<�;�_�z�}�W���Y����R
��[�����;�!�u�;��<�Ϗ�����^��E����4�u�u�;�w�}�6��s���F�N��U���4�0�;�'�:�3�W����Ƹ�VF��Y��ʷ�:�>�=�"�:�>�W�������^����U���u�u�u�u�w�}�����ƪ�AF��T�����4�6�9�!�8�s�Z�ԑT���F�N��9���&��0�3�9�8�1�������pF��DN�����6�0�u�'�:�)�Ͻ�������DחX���u�u�u�u�5�;��������@����U���6��6�:�1����Y������S��U���!�4�u�=�]�p�W���Y�����Q�����u�:�>� �w�<�W����ƭ���E��U���:�:�u�=�w�8����s��ƴF�N��U���&�<�=�&��8��������g��z/�����&�!�0�6�9�/�ϫ��ƥ��������_�x�u�u�w�}�WϽ�����Z���� ���7�u�0�#�4�9��������r%��EN�����:�!�0�;�/�s�Z�ԑT���F�N��6����6�0��9�.��������G�������:�u�4�,�4�>����ӕ��F
��D�����u�u�u�u�w�}��������TF��Q��U���&�;�&�!�2�-�����Ƹ�VF��O��4���u�3�!�<�]�p�W���Y���+����U���<�=�1�4�;�2�W���Y����U��R ��U·�6� �0�!�2�>�������F�N��Uʥ�4�0�<�u�%�<��������{��R������1�-�:��4�:���Y������DN��6���u�u�u�u�w�}����
������^�������=�&�4�0����Ӈ��	��^����� �4�<�;�z�}�W���Y���P��R�X�߇x�u�u�u�w�}��������_��C��ʡ�<�u�9�6�w�5�Ϫ�Y����VF��RN�����;�u�;�u��)�>���T���F�N�����0�u�:�!�2�9��������V�CחX���u�u�u�u�$�8��������]F��[�����u�9�6�u�?�)��������\F��V�����<�2�3�:�w�5�}��Y���F�
��ʸ�8�'�0�{�w�5�Ϭ��ƭ�W��DN��U���'�8�;�0�w�2�W���ӈ����T�����_�x�u�u�w�}�WϪ��ƻ�_
��RN�����,�!�0���W�Z��Y���F�N�����1�'�&��#�)��������V��G�����;�u�;�!� �<�W�������W��D���߇x�u�u�u�w�}����ӑ��[F��EN��ʻ�-�u�:�%�#�)���T���F�N��U����6�8�;�w�3�W�������bF��RN��ʱ�!�u�=�u�6�}��������A	��C�����<� �_�x�w�}�W���YӖ��P��^ �� ���{�u�=�&�3�)�W���ӄ��R��SN��U���u�4�4�6�:�(���� Ӓ��@FǶN��U���u�u� �<�y�p�}��Y���F������ ��9�1�>�9����
ӑ��]F��RN������!�u�;�w���������R
��DN���߇x�u�u�u�w�}��������[��@��U���!�>�;�3�8�}��������A	��D��ʠ�<�u�;�!�2�>����T���F�N�����;�<�4�0� �8�W���Y����_F��C��U���#�9�1�u�$�>�����ƭ�WF��T��:���_�x�u�u�w�}�WϿ�Ӓ�� ��V�����!�1�#�9�2�}��������C��R�����9�6�{�x�]�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���l��^�����0�0�u�:�<�W�W���Y������h�����d�a�4�9�]�}��������F��^�����9�n�u� �2�*��������G��C��1���4�9�_�u�$�}����)����R��X ��1���8�!�'�4�;�W�W�������JF��V�����:� �<�u�$�W�W�������9F������;�=�<�u�w�}�W�������R��N�����3��8�;�#�3����ƥ�G��EG�Uʥ�'�}�u�u�6�8����Y����\	��V �U���&�&�'�0�2�}�MϷ�Y����V��=N��U���%�0�9�u�w�3��������l�N��U���u�&�=�&��>��������]F��D������8�=�&��)�Z�������V�N� ��d�_�u�u��*��������W��X������o�<�u�9�4����H�ƨ�D��^�U��� �g�d�_�w�}�?�������V ��Y
��3���=�&��u�w�3��������W��X����n�u�x�d�y�o�W���
����p��R�����;�u�u�;�"�.����Q�ƨ�D��^�U��� �{�_�u�w�����:����\��YN�����;�_�u�u�w�.����)����e��SN����:�9�4�n�w�}��������@��� ���2�0�}��:�5��������W	��C��\���x� �f�d�]�}�W���
����~��_��:���4�<�u�u�"�}������ƹF��y��8���=�&��!�m�2�ϫ�
����WN��B�����<�&�d�1� �)�W���Y����U�d��U�ߊu�u��!������Cӏ��Q	��R�����u��!���g��������W��S�����|�u�x��o�l�W���
����z��N��U���;�1�d�u�8�3���B���`W��d��Uʦ�0�1�1�'�$��W���ӓ��Z��SF����!�u�|�u�z��G��s���9F������1�0�&� �w�2�ϫ�
����WN��S�����|�u�x� �g�l�}���Y���9F������;�u�u�;�$�:����Nӂ��]��G�U����m�f�u�w�.����0�����D�����b�1�"�!�w�t�W��Y���� l�NךU����6�8� ��1�������\	��V �U���&�6� ��#�>�>������Z��SF�U���;�:�e�n�w�p�$��J�����T�� ���9�u�u� �w�4����M�ƨ�D��^�U���u�a�{�_�w�}�6�������\��B�����1�a�u�:�9�2�G��Y����^�=N��U���6�8� ��m�2�ϭ�����Q��X����|�u�x�u�c�s�}���Y����G"��g�� ���n�_�'�=�#�>����+����UF��V�����:� �<�u�$�}�}���Yӕ��]��D;�����0��%�u�m�?�������G��d�����4�u��&�#�/��������	F��X����u�4�&�n�w�.����Y����G��t��1���,�o��:�2�3��������\��XN�U��}�!�0�&�j�}����P���@��V��6����4�0� ��1��������q	��R�����'�c�1�"�#�}�^��Yۉ��V��
P�����|�_�u�<�9�1��������e��S*�����u�:�9�4��>����Hӂ��]��G��H���!�0�&�h�w�<����s��ƹ��E�����0�%�o�&�%�3�L���s���#��B�����u�=�&�u�>�3�Ϸ�Y����^��R
�����:�=�'�u�%�0����Ӷ��P3��C��ʡ�4�u�=�_�w�p��������V
�������!�u�4�!�>�(�ϵ��ƣ���D������1�0�&�w�4��������A��d��U���u�_�u�x�?�2�(���
����9F��^	��ʦ�4�6�=�&��)�W���������Z-�����&��!�x�w�2����I��ƹ��Y�����6�=�&��#�<�������R��N�����u��0�3�"�g����������Y��E��u�&�2�4�w���������	F��P ��]��1�"�!�u�~�W�W�������w��z�� ���u�<�;�1�f�}�������9F��^	��ʦ�0�!�4��6�8�����ƹ�@��R
��;���=�&��!�z�}�������9F��^	��ʦ�0�!�4��6�8��������_\��X����u�&�2�4�w���������	F��X���ߊu�x�=�:��4����s����]lǻC�6���!�u�=�u�8�)��������F�A������4�!�0��2�"���:����\
ǻC�����
�u��&�6�)��������Gl�C�����4�&�0�!�6���������Z��y��8���=�&��!�6�4�;���Y����[	��h��;����6�=�&��)��������[��x���ߊu�'�6��4�/��������A	��N�����u�:�>��6�)��������G%��C��U��_�u�u�8�)����Q���F��e�����u�u�u�u�w�}�W���Y���F��R��Y���u�u�u�u�w�}�W���Y���K��YN�����4�_�u�u�w�<�������F�N��U���u�u�u�k��0�������F�N��U���u�u�u�x�w�3�W���&����Pl�N�����!�'�u�u�w�}�W���Y���F�
P�� ����&�!�u�w�}�W���Y���F�C����7�:�0�;�w�}�Wϭ�����]��Z��U���u�u�u�u�w�`�W�������P��R ��U���u�u�u�u�w�}�ZϷ�Yӓ��Z��SF�� �ߊu�u�u�� �.�4�������K ��c��8���u�k�&�:�2�)����0����u	��_��4���u�x�u�;�w�3��������Wl�N�����=�&��0�1�3��������~'��
P��=���0�!�:�3��9����-����r%�C���� �&�2�0��l����Y����p��t�����;�&�;�u�w�}�W���D�ƿ�R
��N����� ��0�u�w�}�W���Y����]F��Y�����b�1�_�u�w�}�$�������V0��^
��U���u�u�u�u�i�.����)����e��SB��U���u�u�u�u�z�}��������]l�N�����'��4�0�w�}�W���Y���F�
P��&���!�=�&�y�w�}�W���Y���F�C���� �&�2�0������Y����}��z������!�4�<�w�}�W���D�ƿ�V��V����� ��9�1�4�q�W���Y����F��X���ߊu�u�u��/�����
����F�N��U���u�k�&�0�#�<�'�������P
�N��U���u�x�u� �w�3����ۍ��^l�N�����!�'��9�w�}�W���Y���F�
P��'���4�!�4�6�w�}�W���Y���F�C����7�:�0�;�w�}�Wϭ�����R��B�����u�u�u�u�w�`�W�������@��C8�����u�u�u�u�w�}�Zϱ�ӄ��_��=N��U����9��4�2�(�W���Y���F�N��Kʦ�4�6�=�&��)�L���Y���F�N��X��� �u�;�<�9�9����s����}��z������!�4�<�w�`��������[��x������9�_�u��%�:�������F�
N�����4��4�0�"���ԜY���l�C�����0�!�0�6�2�;����Ӆ��P��C��U���#�:�>�0��<����:����p��=N��X���:�
�u��6�8�ϭ�����R��BךU���6��6�:�1�����Y����G��X��3���!�0��0�1�<����-��ƹF��R �����4�u�_�u�w�}�4�������]��Y��H����0�3�0��.����P����������_�u�u�:�#�0����Y�����D��U���u�h�u��$�)�W���Y���K��YN�����4�_�u�u�w�<�������[�d�����>�u�u�u�z�}��������T��N��Uʦ�&��!�:�1�}�Iϭ�
����p	��QB��U���<�u�7�:�2�3�W���Yӕ��R��YN��U��u��9��6�8���Y����]F��Y�����>� ��9��<����
����\��XN����u�u��0�1�(�W���D�ƿ�\��x��N���u�x�u� �w�4����K�ƨ�D��^��U���u�u�u�u�]�}�Zώ�	����VF��R�����9�u�;�u��1�'�������R
�������0�&�!�u�8�}����Y���P	��Q�����6�9� �4�>�3���� ���C��R�����0�y�4�%�2�1�^�������9F������0�|�!�0�]�}�W���+����A��[�����i�u�:�=�%�}�Iϸ����9F�N��6����4�0� ��1�������N��_��U��3�9�0�n�w�}����Ӕ��Z��R
��]���%�0�9�|�#�8�}���Y�ƿ�V��E�����9�,�i�u��.��������_��D<������9��9�.�5���Y����G	�N�����!�'��9�l�}�W���
����c��R!��#���1�0�4�u�j�.��������F��[�����}��9��6�8��������_��_��X���:�;�:�e�w�}�4���)����|��V��N���u�0�1�<�l�}����	����@��=N��Xʇ�&�4�!�!�2�0����Y����VF��^ ��ʢ�0�u��&�#�9�������F��X��´�0�0�y�4�'�8����Yӄ��ZǻN��´�0�0�|�!�2�W�W���Y����V��^�����&�u�h�3�;�8�}���Y�ƿ�@��R��%���u�h�!� �l�}�Wϻ�
����Z��P1�����4�%�0�9�~�)��ԜY���@3��E<�����%�u�h�&�$�/����B���F��e�����!��1�0�$�a�W�������V��G�����:�u� �0��.��ԜY�Ʃ�WF��d�����%�:�0�&�w�}�W��Y����G��_�����8�8�'�_�w�p�9���Y����4��C��6���u�;�u�4�4�5��������WF��RN�����1�7�u�"�w�1���� ����F��_�����:�0�7�6�"�8��������F������'�4�u�4�?�4�W���Y����XF��T�����!�'�!�4�w�5�W�������V��T�� ���<�;�%�!�y�}�Ϸ�Y����C��C�����_�u�x�!�2�8����
����_��V��ʡ�4�u�0�4�>�:��������VF�������4�!�'�!�2�0����Y����l�C�����0��4�!�2���������w��z���ߊu�x�=�:��}�;���+����W��D��U���&�4�!�4�4�8����P�����X��U���1�!��4��9����
����c��R!��#���1�0�4�}�~�}�Z¨�������V
�����&�;�&�0�3�9����0���K��X��ʦ�4�4� ��$�<����6����F�A�����&�4�4� ��.��������bl�s��8���'�o�0�!�#�}����?����w��V�����,�}��|�w�}����Y����l�N�����0�u�u�u�w�}�W���GӇ��@��N��U���u�u�u�u�w�}�W��Y���Q	��R��U���u��8�9��6�W���Y���X��V�����y�u�u�u�w�}�W���Y���F��N�����2�6�u�u�w�.����.����r��R��H����&�!�'�#�����
���F�N��Xʼ�u�7�:�0�9�}�W���
����a��v
�����;�h�u��$�<��������JN��N��U���u�x�<�u�5�2����Y�����S��'����1�0�&�j�}�4���)����|��V��1���,�d�y�u�z�4�Wϼ�����9F�N��'����1�0�&�9�}�W��Y����W'��E��<���u�u�u�u�w�}�W������]��Y��Lʱ�"�!�u�|�w�}�Wϭ�����e��SN��U���h�u��!������Y���F�N��U���x�<�u�7�8�8����Y����w��~ ��U���u�u�u�h�w�����0���F�N��U���u�u�u�x�>�}����������Y��E�ߊu�u�u��#��&���Y���F�	N�����;�y�u�u�w�}�W���Y���F���U���;�1�d�u�8�3���s���F��V�� ���u�u�u�u�w�c��������F��N��U���u�u�u�u�z�}��������W��S�����|�u�u�u�$�<����(���F�N��U���!��8� ��}�W���Y���F�C����&�2�0�}�`�9� ���Y��ƹF������1�0�&� �w�}�J���+����W��D����u�u�u�u�w�}�Zϱ�ӓ��Z��SF����!�u�|�u�w�}�W���s���%��V��������u�z�+����Ӡ��P��D�����4�u�4��w�p��������a��V�����&�0�!�'��1�3��� ە��@��C-�����4�r�<�=�]�}�Z�������@"��V8������9��4�2�(�!�������JN��V������!�4�<��1�ȶ���ƹK��_��*����0�3�;�$�2���������X��U���!��u��#�����0�����X��U���6�8�;�&�4�(�>���Y����[	��h��4���8� �u��4�0����Y����[	��h��4���8� ��9�$�>��������9F��V��U���<�,�"�'�y�/����
����V��TN��!���u�u�2�;�%�>����Q���F��q�����=�<�u�k�<�4����:����F�N��Uʷ�:�0�;�u�w�-�������F�N������>�u�u�i�����:���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���x�u�;�u�#��W���Yӕ��G��[��U��u��9��6�8��������_��D-�����&��!�4�>���������F�N��Uʷ�:�_�u�u�w���������[�D<������9��9�.�.��������P"��V�����y�u�u�u�w�}�W���Tӏ����[d��U���&�4�4�;�w�}�W���
����~��B��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�x�w�3�W������F��t�����u�u�h�u��8����U���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���<�u�&�2�]�}�W���8����z�N��Kʦ�6� ���w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���K��YN�����u�u�u�&�4�(�8���Y�����T�� ���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�Z����ƿ�TǻN��U���6�8� ��;�`�W�������G*��~G�U���u�u�u�u�w�}�W���Y���F�N��U���u�u�x�:�#�.��ԜY��ƹK�t�����=�u�u��]�}�Z�������u��C<�����0��6��4�W�W�������RF��R�����9�u��&�6�)��������@4��C��6����9�,�=�0�t�W������l��s��#���1�&�4�6�?�.�8�������V
�������4�0� ��;�9����^����l�C�����4�&�:�3��}�4�������F�A�����&�4�4�;�$�<����6����F�A�����&�6� ��w��������K��X��ʦ�6� ��!�$�>�������K��X��ʦ�6� ��!�4�}�6�������P
��N����0�!�!�u�8�6�1�������^��E#��U��_�u�u�2�8�������F�N�������4�;�j�}�1�������R��N�U���u�:�9�4�]�}�W���Ӌ��NǻN��U���%�0�9�u�w�`�W���	����XJ�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�x�<�w�.��ԜY���@"��V8�����u�k�&�4�4�5��������W"��V��6����4�0� ��1��������T�N�U���u�:�9�u�w�}��������R
��
P��'���4�!�4�6�2�<�_���
����p��s��ͽ�2�|�u�u�w�}�W���Y���Z�U�����u�u��!��}�W���D�ƿ�R��R�����u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�p����
����F�N������u�u�u�i�.����6���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���x�u�;�u�>�3�W���Yӕ��P��YN��U��u��6�8�9�q�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��Uʦ�2�_�u�u�w��������[�D/�� ���!�y�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���TӉ����Yd��U���&�6� ��#�>�W���
����^)��{��\���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�x�w�(�W������l�C�����<�0�!�0�$�8����)����|��V��9���&�2�4�u�8�>����Y����F��C8�����u�=�&�6�:�8����
���F��EN��ʶ�0�3�6�0�#�>������������U���u�0�4�{�w�-����
ۇ��@��=�����9�|�u�7�0�3�W����έ�V��N�����u�u�u�&�4�(�8�������V
��R��]���0�&�h�u�6�.�^�ԜY�Ʃ�@��E�����1�0��8�;�������ƹF������ ��9�1�2�<�W��
����^)��a�����4�}��6�:�(�!�������JA��P��U���;�:�e�u�w���������V)��a�����n�u�u�0�3�4�L�������A	��D�U���_�u��6�:�(�!������@'��B�����<��9�,�$�>��������W"��V�����n�u�_�;�w�	�L�