-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����A��s�����9�6��%�!�9�Z�������	F��_ �����8�;�4�1��.�W�������K��E������:�0�!�w����MƴƴF��C�D��� �0�g�d�]�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�=C�]���g�d�u�:�.�4��������R
��Y�� ���!�u�:�%�%�)��ԑTӧ��4��_��'���'�0�_�x��)����Y����A��Y��<���'�4�u�;�8�0����s���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���_�x��'�8�8�Wϊ��ƪ�_��X�����!�&�!�0�'�2�����Ʈ�\��Q�����3�4�!�:�6�W�Z���Y���F��R�����u� �;�;�w�3�ϸ�
����P
��\N��U���u�0�9�&�:�1�W������F�N��U���:�4�;�u��}����Y����R��X �����4�%�0�9�w�2����Yӯ��K�N��U���u�=�;�8�!�.��������G	��_�����9�u�:�4�9�*�����ơ�_��[�����u�u�u�u�w�+����Ӊ��`��[���߇x�u�u�u�w�}�#���	����@��PN��U���0�<�u�=�w�+����Y����Z��Y
�����!�0�:�!�"�W�Z���Y���F��V�����'�;�3�'�2�}�����Ƹ�VF��Z��6���1�8�<�{�z�W�Z���Y���F��x�����>�4�!�'�>�9����
ӎ����NN�����>�6�6�0�w�5�������F�N��U���:�u�4�=��0�������9K�N��U���u�>�;� ��0��������_��Y
�����=�"�8�;�w�<����Y������^��X���u�u�u�u�w�8����
ӏ��G��D*�����z�u�'�4�$�}�3���0�����������x�u�u�u�w�}�W�������R��YN�����9�u�z�u�6�/�W���Ӄ��^�������4�'�,�<�]�p�W���Y�����D�����u�<�3�'�9�}��������P��R@�����=�&�'�4�8�W�Z���Y���F��~ �����%�0��'�.�1�W����Ƹ���D�����!�4�u�'�2�(�Ϫ�s���F�N��U���0�6�:�>�6�)��ԑT���F�N��Uʁ�<�u�:� �2�.����Y�Ƣ�DF��[�����;�0�0�,�#�0�W�������R��V�����u�u�u�u�w�<����
����GF��[�����6�9� �4�2�)�ϸ�����\��BחX���u�u�u�u�$�>�����ɝ�\��B�����<�u�4�<�w�5�ϭ�����F��[�����'�&�u�� �p�W���Y���F��C��ʦ�<�!�1�<�#�}��������A��D��ʷ�u�&�0�!�9�}�3���0����ZǶN��U���u�u�"�!�w�<��������]F��V�����{�x�_�x�w�}�W���YӲ����B�����7�u�0�0�w�4�Ϫ�Ӈ��]��X ��ʴ�#�%�4�0�2�s�Z���Y���F�c�����9�u�4�u�2�/��������JF��D�����&�&�'�0�2�s�Z���Y���F�y��U���u��1�4�%�0�����ơ�@��v������9�1�1�%�3�W���Y����Al�N��U���u�u� �0��.�Ϫ�Y����WF��NN�����&�6� ��#�<���T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���_�<�'�'�w�8��������F��RN�����!�
�:�<��l�C������F��^��[���0�<�
�!�y�1�L�������\��g�����9�!�0��'�<��ԜY����D	��>��1���4�9�_�u�$�}����)����R��X ��1���8�!�'�4�;�W�����Ɗ�R��R�����:�>�:�u�$�}�������F�\'�� ���8�9�&�0��>����ƥ�G��EN��H��_�u�u��2�>��������F�N����;�0�0�u�m�}�^�ԜY����l�N�����4�0�0�u�w�3��������F�d�����>�o�<�u�#�����B���)��E-��U���;�&�1�9�0�>�}���Y����A4��R��U���7�:�0�;�]�}�Wϭ�
����p	��QN����:�9�4�n�w�}����
����A��Y��U��� �&�2�0������
����@K��S�����|�u�x� �d�l�}���Y����P%��[������0�o�<�w�3��������\��XN�N���x�m�m�_�w�}�$�������V0��^
��U���7�:�0�;�]�}�W�������R��N��U���<�;�1�>�"����������Y��E��u�x�g�{�e�W�W���=����]0��^
��U���7�:�0�;�]�}�W�������\��YN�����d��'�,�#�6����*����V��E-�����u�:�;�:�g�f�Z���H����F�D*�����u�u�;��0�8�Fן�������G�����0��'�,�;�p�W������]�N��M��u�u�&�0�3�9����Y�ƥ���^	����1�"�!�u�~�}�Zϋ�I����9F������ ��9�1�m�2�ϼ�����l�N������!�u�u�"�}��������W	��C��\���x�u�a�{�]�}�W�������G7���U���;�1�a�u�8�3���P���F��@�����4�!�0��2�5�������9l��T�����'�u��u�1���������P$��T��ʼ�_�u�x��;�9�>�������G��(�����u�:�u�=�$�0����Y����F��SN�U���0�u�4� �$�5�������K��R�����0�{�u�&�5�$�ϑ�:����P��e�����<�u�;�0�2�}����Y�ƨ�D��\�U���u�0�<�,�<�+��������G	��^��ʧ�;�0�1�3�9�9��������\��V�����2�
�{�u�z�}��������G��B�����u� �%�'�$�.��������9F��X �����>�0�<�,�!�1�1�������|��\(�����4�2�
�_�w�}�W���Y���F�N��U���u�u�o�u�!�1�1�������T�������:�>�4�!�%�f�}���TӰ��Z��B��ʺ�u�4�%�0�w�8�W����ƪ�AF��^�����0�4�0�d�#�}�8�������u��X�:���'�u�x�u�6�(�Ͻ�����Q��E�����:�4�&�;�;�}�%�������V��P�Uʦ�7�,�0��4�<����Y����]��R�����u��0�6�8�6����ӂ��]��UךU����'�3�u��-����	����V��T�����;�'�;�0�3�;�����Ɵ�P4��P��[���6�;�!�;�w�����0����`��N�����;�0�!�u�w�}�W���Y���F�N��U���o�u�%��9�8�ǵ�����R��R�����9�|�_�u�z�}��������	��C�����:�<�2�!�8�+����
ӑ����R�����0�0�!�1�]�}�Zϱ�����`����U���0�6�:�>�6�)����HӠ����������;�u�4�]�}�Zϵ�����\��V��ʓ�&�u�:�0�3�)��������V��^��U���!�0�%�:�2�.�W��Y������DN�����<�;�9�{�w�.����Y����R/��N ��Oʗ�:�0�;�0�#�/��������X ��C�����!�u�|�o�w�2����Y����R
��UךU���;�9�:� �'�)����CӤ��_��a������0�6�:�<�<����Hӂ��]��G��H���!�0�&�h�w�<����s����Z��[N�����0�0��%�w�}����������RUװUʦ�2�4�u��6�8��������Z��N�����0�}��8�?�.�5���T�ƨ�D��^��O���:�=�'�u�i�z�P��Y�˙� H��=N�����9�&�4�6�.�1��������c��T�����;�1�b�1� �)�W���C����G��DN��U��|�u�x� �y�W�W�������`��C>�����9�1�<�0�m�?�������U��RUךU���;�9�&�!�%����������^	��¾� ��4�0�>�.�FϺ�����O�
N�����&�h�u�e�~�}�Z�J����F��P ��U���!���9�3�4�������R�
N�����_�u�<�;�;�.��������zF��d�����'�,�!�<�3��������c��N��X���:�;�:�e�w�`�_������F��C����r�r�|�u�z��O��Yӕ��]��D*�����<�0�u�u�>�3��������GN��Y��&���9�&�0��4�8�FϺ�����O�
N�����&�h�u�:�?�/�W���I���K�d_�D���&�2�4�u��<�6�������C������1�l�1�"�#�}�^��Yۉ��V��
P��E���u�x� �e�f�W�W�������f��[�����<�0�o�7�8�8���Y����V]ǑN�����u� �0��$�)�Mϼ�����\�C��N�ߊu�<�;�9�8�5��������]������1�>� ��6�8����Hӂ��]��G��H���!�0�&�h�w�m�^���T޳��W��N�����u��9��4�8�:���
����	F��D�����u�:�;�:�g�}�J�������[�^��N���x�m�m�u�$�:����*����c��R8�����u�:�9�4�w�`�������@��V��&���!�=�&�u�w�3����ۍ��^6��D�����u�:�;�:�g�}�J�������[�^��N���x�g�{�g�w�.����Y����R/��V��U���:�9�4�u�j�;����s�ƿ�T��������9�1�4�2�}������ƓF��P ��U���!���o��:���8����l��~ �����%�0��'�.�1�Z�������V�S�����'�u�k�}�#�8���^���F�=�[�ߊu�<�;�9�8�<����Y�Ɵ�T��V�����!�>�;� ��0��������_�
�����e�u�h�}�#�8���Yۉ��V��
P��R���u�x��m�f�}�����ƣ�R��Y=�����u�u�<�;�3�u�@Ϻ�����O��N�����u��!���/����Cӕ��]��_����!�u�|�_�w�4��������r��R��Oʠ�&�2�0�}�w�2����I����N��_��U��r�r�n�x�w�l�Y��Yӕ��]��X;��4���:�3�u�u�8�1����DӀ��@��=N�����9�:�6� ��)����)����	F��X����u�4�&�n�w�.����Y����F��C>�����u�<�;�1�c�}�������	[�X�����k�r�r�n�z�}�C���s�ƿ�T������� ��%��m�.����Q����\��XN�U��}�!�0�&�j�}�G���Y����S�=d�����4�u��6�:�(�!�������	F��S1�����o�u�e�n�w�.����Y����F��C"��<��&�2�0�}�c�9� ���Y���F��C����u�e�|�u�z��B��Yӕ��]��D/�� ���!�6��o�$�:����Mӂ��]��G��H���!�0�&�h�w�m�^���Tӵ��VǑN�����u��4�9�w�}��������G	��N�����u�|�_�u�$�:����=����]/��R� ���2�0�}�:�e�8����6����_	��q�����:�;�:�e�l�}�����ƣ�J��X��Oʠ�&�2�0�}�8�o����Q����A��T�����|�:�;�:�g�f�Wϭ�����@#��U�� ���!��u�:�;�<�L�ԜY�˺�\	��D�����_�u�<�;�;�2����6������Y��A���:�;�:�e�l�}�����ƣ�P��x��Oʦ�2�0�}�a�3�*����P���@��V��4���8� ��9�3�}������ƹ��Y�����6�:�;��;�9�W�������9F������<�0�1�_�w�)�����Ƨ�V������_�u�x�u�?�.�W�������R��VN�����u�!�'�7�#�}�ϻ�
����G����ʱ�;�!�2�!�w�p�W�������]��d<��G���u�=�'�u�2�9�W����ƭ�]	��X	��U���=�7�!�0�9�)����T�Ɵ�^��t������0��>�3�0��������Z��P@ךU���'�7�!�u�2�-����,����V��N�����u�&�w�'�2�f�WϿ�����G��R������4�0�;�%�0���
����_F��L�� ���_�u�!�'�5�)�W���	Ӊ��\%��T-�����<� ��0�w�4��������A��d�����<� �0�>�2�}�ϱ�����[��N�����u�&�w�'�2�f�WϿ�����G��R������!���w�4��������A��d�����<� �0�>�2�}�ϱ�����b\��^	��ʼ�u�!� �w�]�}��������X�������1�1�'�&�m�.����Y���G��UךU���'�7�!�u�2�-����,����G%��Q����4�u�&�w�%�8�L�������Q����ʺ�u��4�!�?�.�!����ƿ�T����W���0�n�u�4�#�4��������\ ��s��<���9�1�u�<�9�1��������lǻC�!���0�&�2�4�w�<�Ͽ�[����F��C�� ���!�u�;� �2�)��������\��	�����x�&�6�0�w�3�ύ�5�Կ�F��R�����&�!�u�0�6�3�W����Ƽ�G��R�����=�_�u�x��8�4�������R��R-��U���4�;�u�:�w�4����s�ƭ�G��B�����u�3�&�6�"���������	F��P ��U���w�'�0�n�w�<��������V��X��4���8� ��9�m�.����Y���G��UךU���'�7�!�u�2�-����8����|��T��U���;�9�<�u�#�(�U�ԶY���v��E�����!�0�&�;�w�4����ӕ��]��S�����0�u�8�9�:�3��������a*��Q�����;�_�u�!�%�?��������UF��V�����6�u�<�;�;�4�Wͪ�����F��C�� ���>�0�u�3�8�(���� ����@��V�����'�0�n�_�2�4�}���TӪ��P��_�����u�<�;�9�w�3����*����V%��
�����7�3�'�u�?�$����
����G	ǻC�����0��>�3�0���Y������S��U���0�&�'�u�?�/�W���ӈ��_	��Td��X���4�=�7�!�2�3��������]��X�����2�u��!�w�5�Ϫ�����Z��[�����4�0�_�u�z�?�W�������VF��P ��U���!�1�0�u�8�}����ӓ��Z
��R�����,�9�&�4�#�/����	����@��N�U���4�&�'�&�w�	��������@F��V�����:�u�=�u�9�(�W���Y����_��B��ʡ�0�'�&�!�w�p�W�������9F��E�������2��$�)�$�������l�U�����u�<�}���:�%����Ƹ�VǻN��U���4�9�u�h��)����D�ƪ�_��d��U���&�&�'�0�2�����DӒ��V]ǻN��U���4�!�=�&��1������� ��D�U���u�&�4�4�9�<����	��� ��D�U���u�&�=�&��>��������Z������h�u�e�|�]�}�W���:����J��D#�� ���0�<�0�i�w�2����Y���A�=N��U����4�!�=�$�����D�Σ�[��S�R��n�u�u�u�$�<��������[�X�����k�}�!�0�$�`�W��P��ƹF�������%��i�w�2����Y���\��E��K��r�|�_�u�w�}�%���8����@��G��H���!�0�&�h�w�m�^�ԜY���@3��v������%�u�h�1�1��ԜY�Ʃ�@��E�����1�0��8�;�������ƹF������u�h�&�;�5�8��������Z��N�����u�|�s�!�"�f�W���Yӏ��@#��U�����7�0�=�2�~�}����Y���F��b��'���!�<�0�i�w�����
����F�N�����'��4�0�6�4�'���Y���@5��E�����4�<�n�u�w�}�Wϭ�����e��S>����u��!���1��ԜY���F��_��<���0�0�!�<�2�a�W�������P��R �����u�u�u��;�����4����|��^��I����9��6�2�������ƹF�N��&���!�=�&��'�}�Jϭ�����[��d��U���u�&�4�4�9�4����Dӕ��G��~UךU���u�u��!������E�ƿ�R��Y?�U���u�u�&�0�3�9����)����[��e��4���0�&�_�u�w�}�W�������\��g��U��&�&��!�8�;�L���Y����]��QUךU���;�u�3�_�w�3�W�������9l�C�����u�=�u�;�"�}�����ƥ���!�����u�:�4�;�w�	����
ӂ��VF���� ���u�x�u�=�%�}�Ͽ��ˠ�T��G��U���"�0�u�=�w�2��������Z��P@ךU���6�&�}���:�%���ߩ��A%��d�����;�u�u�<���1���+����F��R ךU���u� �0��$�)�K�������F�N������4�0�4�>�}�Jϸ�����F�N������6�0�0�#�a�WǱ�����X�I����u�u��9��>��������VF�F�����u�k�r�r�l�}�W�������G6��D��H���!�0�&�h�w�m�^�ԜY���\"��V'�����u�h�3�9�2�W�W���Y����R/��R��]���0�&�h�u�8�5����G����O��N��Uʺ�4�4�;�u�j�u����
���	��R��H���e�|�n�u�w�}��������V��S�����'�u�k�r�p�f�W���YӉ��V'��t����u�4�&�n�w�}����Ӕ��Z��R
��]���'�9�|�!�2�W�W���Y����A4��R��Hʦ�&�'�0�0��-�L���Y����`��C>�����9�1�i�u�$�)��������_��^�����u�u��4�2�3���������V�����8�;��%�l�}�W�������p��R�����;�u�h�&�6�>����
����@)��g��N���u�u�:�!�%�����E�ƿ�G��g�����0�_�u�u�w�����/����Z�D*�����4�<��%�l�}�W�������z��S��1�����%��]�}�W���=����]7�
N�����;�<�0�n�w�}�Wϱ�����W��DN�U���4��1�0�$�4��ԜY���\3��v�����u�h�&�&��)����)����9F���U���_�u�;�u�%�>���s���%��V�����:�4�4�;�.�>�����Ƹ�R��R��U���u�#�'�9�w��W���Ӓ��@��[ךU���1�!�u�'�:�)�ύ�����_��X������0�!�u�?�}�8�������PF��P ��U���!�!�9�&�w�p�W���Y����p
��X�� ����u�=�;�#�}����Y����W�������u�=�u� �'�)�$�������9F�N�����u��u�0�w�)��������l�C�����0��0�6�8�6��������]��=N��X���:�
�u��2�>����������R�����4�!�'�u�z�+����Ӎ��F��V�����u�f�w�u�z�+����Ӈ��@��V"�����0�0�_�u�z�5����Y����p
��d�����>�u�x�#�8�6�ϱ�����\5��T-���ߊu�x�=�:��}�4�������WF��N ������9�1�u�z�+����Ӊ��@��\+�����!�:�0�_�w�+��������`��t�����o�0�!�!�w�2��������P��P=�����;�0�u���W�W�������PF��GN��U���u�>�#�'�;�>�1��������R�����4�!�'�u�z�}��������AF��]ךU���u�� �!�6�����Y���U��N��U���u�u�u�u�z�4�Wϭ�����	[�^��U���%�'�u�4�w�W�W���Y����V�N��U���u�k�4�#�'�<����U���K�^ �����0�;�u�u�w��������F�N��U���%�0�9�y�w�}�W���Tӏ����h���ߊu�u�u�#�%�1�W���Y���[�x��6���u�u�u�u�w�p�W���Y����_	��Td��U���:�:�;�u�w�}�W���Y����`��t�����u�u�u�x�8�)��������_	��[��D¾�#�'�9�6��>�������F��t�����<�u�u�u�j�}�$���:����e��SB��X��� �u�:�9�6�W�W���Y����V%��r
��;���u�k�:�0�~�}�W���Y���K�X�����0�;�_�u�z������Ƹ�VF��Y�����9�u�:�8�<�}����Ӄ��Z��C�����u��!���3�W���	����Z��=N��Xʾ�#�'�9�6��>����Y�Ư�P
��N�� ���!�,�6�>�!�/����?����AF��T��[���x�u�:�0�#�<�W�������]��DN��ʦ�;�0�u�:�#�8�$���������RN�����4�0�,�4�#�/����	����@��=N��Xʁ�0�0�:�0� �}����*����\��a��ʡ�u�4�>�4�.�(�����ƣ�J��X��U���%�'�&�;�y�}����������P������0��>�]�}����s���Z ��{�����&�!�u�=�9�}�W�������z��Y��I���:�=�'�u�i�;����B���F��s��<���1�-�u�h��)����D���O��N��Uʺ� �%�!�,�4�a�WǱ�����X��V��\�ߊu�u�9�<�w�4��������|��t��U���;�u�u�u�z�}��������Z��CN�����&�4�0�'�0�.����Y����GF����U���%�0�9�u�8�<����Y���F��SN�����;�!�0��2��Ϻ�����2��DN������0��>�$�:��������T��N��U���u�=�<�u�2�}����
Ӊ��G��D�����1�0�:�u�!�/��������RF��D�����u�u�x�0�0�}�ύ�����_��Y
�����!�0�'�#�;�8��������X ��C�����0�{�u�u�w�p�W���Y����Z��=��U���u� �0�u�9�2�ϭ�����@��V�����u��;��"�)�������F�C�����u�;�u��#��$���Y����A��R �����,�9�&�!�w�/����0����`��[�����6�0�u�u�w�p�W���Ӓ��"��VN�����{�u�u�u�z�}�Ͽ�����A	��D��ʰ�6�u�<�;�;�0��������]��@�����:�4�4�;�6�4�W������F�N�����;�,�6�u�w�}�Z���Ӄ��F��C��&���9��>�1�:�4�W���
Ӄ��[F��[����� �u�'�8�#�8��������\ǻN��U���"�u�4�0�#�8�����ƿ�T��DN������!� ��9�s�W���Y���F�N�U���0�<�u�u�>�:����ӏ��F��V�����!�0��;�w�4����Y����R��P ��U���;�u�u�u�z�}�8�������u��X����_�u�u�u�z�}�W���Y���F�N��*���
�u�u�u�w�}�(���&����F�N��U���
�
�
�u�w�}�Z���*����V%��N��*���u�u�u�u���(������F�K1��*���
�u�u�u�w�!�(���&��ƹF�C�U���u�u�u�u�w�}�W���Y�Ɠ�F�h1��Uʊ�u�u�
�u�w��W���&���9��N��*���u�u�x�u��8�4���Y���l9����	���
�)�u�
�+�}�(���Y����F��h��	���u�)�
�u�+��W���Y���F�N��U���u�u�u�
���(���&����l9��h1��*���
�
�
�
���(���&����l9��=N��U���x�u��;��)����&��ƹF�C�U���u�x�u�:�.�>����Y���OF�N��U���)�u�u�)�w�}����YӚ�F��N�U���d�u�u�g�w�}�W��Y���F�N��U���u�u�u�u���W���Y���F�h1��*���u�u�u�u�w��(���Y���K�������;�}�|�f��4���Y����l9��h1��*���u�u�u�
���(���&���F��h1�����u�u�x�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�Wρ�&���F�N��U���
�
�_�u�w�}�Z���=����]5��TF�����d���
���(���&����OF�N��*���
�
�
�)�w�}����&���F�CךU���u�x�u�u�w�}�W���Y���F�N��*���
�
�
�u�w�}�(���&����l9�N��U���
�
�
�
�]�}�W���T�ƣ�R��Y=����u�u��
�w�}�W���Y�ư�l9��KN��U���u�u�)�
��!�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��*���
�
�
�
�w�}�Wρ�&����l9��=N��U���x�u��!���������F��t1��*���
�
�
�
��}�W���Y���O9��h1��U���u�x�_�u�w�}�Z���Y���F�N��Uʊ�
�
�
�
���(���Y���K�������9�1�
�+�}�W���Y���F���*���
�
�
�
���(���&����l9��h1�����u�u�x�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�Wρ�&����l9��h1��*�ߊu�u�u�x�w�����/����9��h1��*���
�
�
�
���(���Y���F�N��U���)�
�
�
���}���Y���9F�N��X����!���;�9����Y���K�N��U���u�u�u�u�w�}�W���Y���F�N��U���
�
�
�u�w�}�Z���Y���F�_��%���
�
�
�
���(���&����l�N��*���
�
�
�
���(���&��ƹF�C�U���u�u�u�u�w�}�W���Y���F�N��U���u�u�
�
���(���Y���K�N��U���u�u�u����(���&����l9��h1��*���u�u�u�u�w�}�(���&����l9��h1�����u�u�x�u�w�}�Z���S���L�D��_�������}�w�]���S���L�D��_�������}�w�]���S��ƹF�C�U���u�u�u�u�w�}�W���&���F�N��Uʊ�
�
�u�u�w�}�W���&����9F�N��X����!� ��9�u�^���Y����l9��h1��*���u�u�u�
���(���&���F��h1��*���
�_�u�u�w�p�W���Y���F�N��U���u�u�u�u���(���Y���F�1��*���u�u�u�u�w�}�(���s���F�N�� ���!�,�6�=�0�t�(���&����OF�N��*���
�
�
�)�w�}����&����l9��=N��U���x�u�u�u�w�}�W���Y���F�N��Uʊ�
�
�u�u�w�p�Wϱ�����F��[��U���u�
�
�
�+�}�WϢ�&����l9��h1��*���
�
�
�
���(���&���F�N��U���u�u�u�u�w�}�W���Y���F�N��*���
�
�
�
���(���Y���F��v������9�1�<�2��(���&����l9��N��U���u�u�u�u�w��(���&����l9��h1ךU���u�x�u�u�w�}�W���Y���l9��h1��U���u�u�u�
���(���Y���F��h1��*���u�u�u�x�w�����:���F��KN��U���u�
�
�
��!�W���Y�ư�l9��h1��U���u�u�)�
���(�ԜY���\"��V'�����i�u��!������=����]5��TI�����u�:�;�:�g�W�W���Y���F�N��U����;�� �#�<��������`��t����>�;� ��:�1����:����O��N��Uʺ�4�4�;�;�2�}�Jϱ� ����F��=N��U����!� ��9�}�Jϱ�����`��������;�r�<�?�l��������9F�N��U���u�u�u�u�w�u�$���:����e��SN��ʺ�,�6�:�;�w�}�8�������u��X��U���_�u�u�;�w�;�}����Ƽ�\��DUװU���u�4�0�!�2�>����ӕ��]����ʺ�4�4�;�,�4�.�W�������D�������u�0�u�4�"�.�W��Y������=�����9�u�:�4�9�}�����ƨ�]A��_��U���2�!�u��6�)����ӄ��R��=N��Xʡ�0��:� �>�����ӑ��_F��Y��U���8�'�u�=�9�)��������@J��Q��U���<�u�&�0�#�9�}���T�΅���[N�����u�!� �!�;�4�Ͻ�����G�������&�0�{�_�w�����/����t��R�����4�;�4�<�w�3�W�������J��X*�����,�6�=�2�~�W�W��Y����\
��V�����8�9�<�9�w�1����
ӏ��@"��V'��Z���;�:�4�&�9�1�W������f��N�U���<�0�<�0�w�8����Y����`��t��ʡ�u�:�!�:�w�5�ϓ�!���K��X�����u��!��������ƿ�R
��EN�����=�u�4�<�"�}�$���:����F��\�� ���u�x�u�=�w�(�W����ƿ�_��DN��U���8�;�u� �w�;������ƹ	��C��&���4��u�i�w�����0ە��_
�������4�%�0��%�$���Y�ƣ�R��Y'�����n�u�:�4�6�3�������[��s��<���&�4�9�'�<�3��������c��N��X���u��!���9����s���%��V�����%�:�0�&�9�}����s���E��\1��3���!�0��:��2����Tސ��\�������4�#�%�4�2�8�}���T����X9��D;�����0�u� �0��.����Tސ��\��=�����9�u�#�'�;�W�W�������RF��D�����3�u� �0�;�����Y����[	��h��%���0�;�'�8�9�}�'�������V��Cd��Xǣ�:�>�4�&�6�>����
����@)�������6�0��;�$�3�}���T����X9��D=�����4�0�4�<�w���������R
��=N��X���:�
�u��6�)����Y����A��V��U���#�:�>�4�$�<��������\"��V'������!�_�u�z�5����Y����R/��������'�4��w�p��������w��~ �����4�;�0�<�;�W�W�������RF��R�����&��u��6�����
�����X��U���6�8� ��;�9��������e��Sd��Xǣ�:�>�4�&�4�(�8���Y����F��C'ךU���=�:�
�u��>����(Ӊ��P��B��Uʓ�4�!�0��8�����CӃ��Z��@��[���6��6�'�4�1����+���F�G��U���u�_�u�u�w�����Y���F�N��H�����2��$�)�W���Y���K��YN�����4�_�u�u�w�����
���F�N��H��� �0��&�#�}�W���Y���K��YN�����4�_�u�u�w�<�������F�N��H���#�'�9�y�w�}�W���Y���K��YN�����:�<�_�u�w�}�"�������U �N��U��u� �0�9��8����Y���F���U���9�4�_�u�w�}�'�������V��CN��U��u��4�0�9�/����U���F���U���<�;�1�>�"����������Y��U���u�&�4�6�.�1��������[�X-�����9�&�<� ��8�W��Y���F��P ��]���:�;�:�e�]�}�W���*����c��R8�����u�h�u��6�)����/����F�N�U���u�:�9�4�]�}�W���*����c��RN��U���u�h�u��6�)����U���F�N�U���u�;�<�;�3�6��������G�
�����u�u�u�&�6�<�������F�S����4�;�4�<��)�[���Y���Z�U�����u�u�u�&�6�<����Y���F�S����4�;�0�<�;�q�W���Y���Z�D�����b�1�"�!�w�t�W���Yӕ��G��fN��U���u�u�u�k�8�<��������bJ�N��U���<�u�&�2�2�u�@Ϻ�����OǻN��U���4��1�0�$�3�W���Y����a��v
�����u�u�u�u�w�p��������]��N�����u�|�u�u�w�.����6����_��N��U��:�6� ��#�<���Y���K�X�����0�;�u�u�w�.����6����F�N��U��:�6� ��#�q�W���Y���K�X�����0�}�a�1� �)�W���Y�����T�� ���u�u�u�u�w�c��������bO��N��U���u�x�:�!�$�:����Mӂ��]��GװU���u�4�6�u�?�}�����ƪ�\��_�����9�u�:�4�9�.�W���Ӓ��JF��RN�����0�u�:�'�4�1�}���Tӏ��G��d�����>�1�8�<�y�}����������P������0��>�]�}����s���Z ��{�����&�!�u�=�9�}�W�������^)��a�����0�i�u�4�$�f�W���YӉ��P��B�����i�u�:�=�%�}�I���^��ƹF������ ��%��k�}�������A��UךU���9�<�u�<�>�:����Q����p
�������u�u�x�u�$�8�ϱ�����F��[�����<�u��6�:�(�!���Ӈ��V����ʼ�u�=�_�u�w�}�ZϪ�����_	�������<�1�"�!�6�}�����Ƹ�VF��Z��6���!�8�;�_�w�}�W�������F��Y��:��� ��;�r�>�5�^Ϫ����F�N������!�4�<��-�W������^)��a���ߊu�u�u�9�2�}�W���YӉ��P��B�����<�0�i�u��>����/����c������� ��!�4�>�f�W���YӃ����=N��U���x��!�=�#�8����Y����F��V �����u��6�8�"���������GǻN��U���:�6� ��#�<��������F�N����� ��!�<�2�}�Jϱ�����F��=N��U���u��6�8�"�����E�ƣ�P��x��N���u�u�0�1�>�f�W�������U]ǻ��U���6�&�n�_�w�p�#���Ӡ����
�����1�1�'�;�w�3�W����Ƹ�VF��D�����:�u��&�#�W�W��8�ƭ�@��^������&�!�8�.�>��������G��[��U���!�<�u�:�"�8�W��Y����VF��Z�����;�;�&�6�9�2�W�������N��gZ��Yʗ�:�>�4�{�2�>�^�ԜY����VF�� ��U���!�!�<�u�2�<��������G	��V�����"�,�!�u�?�}�!Ϙ�>���K��^�����u�:�u�0�3�.��������Z��(��U���!�<�u�:�"�8����ӑ��R��N�U���0�!�4�u�;�}�Ϫ�Ӌ��R��U�����4�u�0�!�2�s�W���Y����Q
��Pd��X��� �4�<�;�6�)�Ͽ�����Z��RC�����0�u�&�6�9�/����Y����[��aN�����8�_�u�x��}����Y����VF�������&�9�;�u�$�)�ύ�����_��^�����1�9�,�u�z�}�����Ƹ�Z��X
���ߊu�x��!�m��W�������G0��^
��ʼ�u�<�4�9�3�u����ӕ��V��D��U���9�u�!�u�z�}�W���Y����A����ʼ�u�<�9�&�6�}����������R�����1�4�&�'�$�W�W��Y���2��"��3���u�<�2�4�w�5��������G����ʃ�9�1�1�'�9�}����s���F�N�����0�%�<�u�6�6�ϸ�Ӈ��_��CN��ʶ�6�0�4�!�%�)�Ϙ�Y����]��R
�Uʦ�;�7�0� �'�)�1��Y����@3��E<����_�u�x�=�8��W�������)��a�����%�u�x�#�8�6�ϵ�����R
�IךU���=�:�
�u��.�Ͽ�����a��Cd��Xǣ�:�>�4�6�9�.��������F��=N��X���:�
�u�9�w�<�������K��X��ʶ�u�:�&�1�8�4�_�������G0��^
�����u�x�#�:�<�<����8����|��V��9���u��!�4�>��������JF��E��3����%�}�!�~�}�WϹ�������FךU���u��&�!�6�}�I���^���F��N�����2�6�o�u�g�W�W�������R�=N��U����&�!�h�w��1���+����F�N��U���u�u�u�u�w�p�W���Y����V��N��Uʶ�;�u�u�k�$�3��������u �N��U���u�u�u�u�w�p��������RǻN��U���u�u�h�u�6�-����U���F�N��U���u�u�u�u�z�}��������T��N��Uʶ�u�u�u�k�#���������r��Z!��#���1�<�0�y�w�p����
����\��=N��U����u�u�h�w���������Z��[G�U���u�u�u�u�w�p�W���Y����_	��TN�U���&�!�4�_�w�p�W�������[��^ ��U���_�u�0�0�6�8��������u ��=N�����u�;�e�!�w���������zA��P�����4�0�u�u�z�+����Ӣ��\��GN������!��:��}�W������l��e�����u�e�_�u�w�p����&�ƭ�V����3����&�!�u�w�p��������v��r �����!� ��_�w�}�Z�������p
��d�����>�u�u�x�!�2�����ƣ�P��x�����}�|�u�u�z�+����Ӆ��@'��B������<�_�u�w�(��������\�������"�'�{��8�������ƹF�	�����u�4�u�_�w�}�W���+����e��
P��E���u�x�<�u�$�9�������V�N��Uʥ�'�u�4�u�]�}�W���Y����V�	N�����4�0�0�y�w�}�W��Y���Q	��R��U���u�u�6�;�w�}�Iϭ�����|��B��Y���u�x�<�u�5�2����Y���F��[��U��u�4�%�0�;�q�W���Y���K��YN�����:�<�_�u�w�}�W���Y���F��T��:���<�0�}�|�w�p�W���Y����_	��Td��U���u�6�u�u�w�c������������N���x�:�!�&�3�1����C�Ƨ�V��a�����u�x�=�:��}�1���=����F��C*�����%�_�u�u�z�5����Y����V��[N��R���u�x�#�:�<�<�����ƭ�E ��V<���ߊu�u�x�=�8��W���Y����Q
��B�����u�u�x�#�8�6�ϝ�ӵ��C
��[ךU���x�=�:�
�w���������c��fF�����u�x�=�:��}�&ϭ�����F��[?��\���u��!� ��)�1���(�Ʃ�G����đ�9�%�&�u�%�1�}���Y�ƫ�]��TN�����u�u�u�u�<�8�������V�N�U���u�!�
�:�>�}�J���^���F��X�����}�u�u�u�w�<����Y������P�����u�u�u�u�z�4�Wϼ�����9F�N��U���u�u�h�u��<��������uJ�N�U���u�:�9�4�]�}�W���Y����F�	N������>�u�u�w�}�W��Y���@��[�����u�u�u�6�w�}�W�������^)��g��$¼�y�u�x�<�w�.������ƹF�N��$���u�h�u��4�0�����Υ�]�C�� ���!�
�:�<�w�`��������9F��Y
�����4�0��;�%�)�8�������R ��dךU����&�2�u�?�}����Y����F��N������!�4�<�w�`��������]N��T��:���4�<��9�l�}��������zF������ ��9�n�w�.����6����[��v������9�n�0�3��;��