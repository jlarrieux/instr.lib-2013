-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����B+�����߇x��!�:�m��Ϝ���ƴF��^	�����'�?�6�o���(��L���"��RT��Gʑ�6�8�0�u�g�l�Z�ԑT���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���6�u�e�d��-����Ө��Z	��[N�����8�;�&��%�2�������r
��e�����0�0�#�1�z�}��������]��B�����;�0�;�9��;������ƴK�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���_�x�x�u�"�-���-����P	��X ��ʼ�%�0�0�!�w�}����	����P��B�����:�7�u�&�3�4�W���T���u/��Q�����<�=�f�u�!�/�������2��DN�����0�!�<�6�"�8�W���Y����U��R ��X���u�0�:�,��2�W�������F��RN�����0�:�,�}�8�}�W���ӑ��W���U���u��a�{�z�W�Zϒ�������-�����<�;�&�_�z�}�#���Y����\��CN�����u�u�:�3�>�4��������_�'�����-�0�!�1�#�<�W���s�����_�����9�6�8�:�2�)� ���Y����A�������<�;�u�4�"�}�ϭ�����]JǶN�����1�&�'�1�;�>����Y����p	��v
��Yʴ�1�!�2�9�w�5�W�������_�����߇x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��s����A�����ߊu�&�u�0�2�.��������P��V�����&�u�0�0�9�0����
����_
��=C����=�&�&�!�6�.��������Z��E�����-�:�0�<�l�1���� ӳ��`/��=��U������:�'�3����8����K��N �����u�'�;�9�#���Զ����JF��z��ʼ�u�_�0�0�>�u�Wϵ�����]%��^ ��U���;�7�:�0�9�g�W���
���9��CFךU���%�0�9�f�w�}�W���ӕ��l
��^����&�:�3�1�%�}�W���Y����G��X	��*���!�'�d�1� �)�W���s�ƿ�p	��`��U���u�o�<�u�#�����B����@%��Q*�����u�u�u�;�$�9��������G	��Y�����:�e�n�u�$���������@F������9�2�6�_�w�.�3���0���F�T��ʦ�1�9�2�6�!�>����Nӂ��]��G�Uʦ��!��!�w�}�W������G��X	��*���!�'�d�u�8�3���B����@"��V8�����u�u�u�;�$�9�������@��C����� �u�o�:�#�.��������F��s��"���u�u�u�o�>�}��������9F��D*����� �u�u�u�w�(�W���&����P]ǻ�����&��u�u�w�}�ϭ�����Z��R����1�"�!�u�~�W�W�������@)��N��Oʺ�!�&�1�9�0�>��������W	��C��\�ߊu�&�6� ��}�W���Y�ƥ���h�����0�!�'�a�w�2����I��ƹ��T��:���u�u�u�u�"�}��������E��X��Bʱ�"�!�u�|�]�}��������Z��CN����&�1�9�2�4�t�}���Y����PU��=d�����!�6� �0����������KF��=d��Xǣ�:�>�&�2�#�/�}���T����X9��P���ߊu�<�;�9�$��������F�N�����2�6�#�6�8�u�W������F��F�����h�r�r�n�]�}����ӕ��R��R!��9���u�o�&�1�;�:���Y���9F��^	��ʦ��1�0�&�"�����Y����_	��T1�����}�u�:�;�8�m�W��Q����A�^��N���&�2�4�u�$�<����*���F���*���<�
�0�!�%�l�W������F��F�����h�r�r�n�w�.����Y����V ��s��U���u�u�!�
�8�4�(������F��@ ��U���o�u�:�=�%�`�P���B����Z��[N��"���0�;�:�7�w�}�W���&����PF��I�N���&�2�4�u�$�<��������F���*���<�
�0�!�%�j��������\������k�e�|�_�5�:��ԜY���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�U���u�&�4�4�6�4�>�ԜY��ƹK���U���!�0�%�4�w�2�W���Ӑ��Z�'�����<�%�!�1�#�}����Y����WJ��_��U���u�:�r�u�%�)�W����Ƹ�VF��C�����,�4�1�=�;�}����*�Ʈ�\��N��R���>�!�_�u�z�1�Ϫ�Ӆ��U ��^��ʾ�0�u�:�9�9�q����Ӓ��JF��G��U���'�u�4�%�2�1�Y���T���K��^ ��U���u�4�4�=�$�<�CϽ�����V
�������u�=�u�$�6�<���� �ƨ�_��N�U���u�4�4�#�;�9�����Ư�P
��C����� �u�<�=�6�}����
����UF��S�����x�"�'�&�w�	�ϸ�����r%��[�����,�u�4�4�!�1�ϼ�Y�Ư�P
��N��ʡ�0�'�&�_�w�p�����Ɓ�p��NN�����u�,�9�{�w�5�ϩ�����F��E�����"�0�u�:�w�2����T�ƭ�����ʺ�u�=�u�<�9�1�W���Ӓ����^ ��ʘ��{�u�x�]�}�Zύ�Y����]��GN�����=�&�6�4�9�2�W�������_��D�����u�=�!�4�2�<�������F��C�����=�<�u�3�$���������@H�c��U���<�%�'�4�#�?����Ӊ��G��=N��Xʣ�'�:�&�%�6�8�W���Y����_���� ���&�8�u�;�#�8�3���A�ƿ�^��B�����_�u�x�4�3�$�ϰ��Ƹ���V��U���u��&�"�2�}��������\�������u�&�r�u�w�p�W������u	��C��U���&�;��0�'�.�Ϫ�Ӆ��P��Y�����;�!�0�<�3�+����s��� ��DN�����u�=�u��c�q��������VF��B�����0�9�u�<�2�4�Ϫ�����@F��[�U���u�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�W��Y���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�=N��Xʑ�!�u�0�:�.�}�Z���T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���KǑN�U���u�4�4�8�:�/�Y�������G	��_�����8�8�'�u�?�3����Y������A��ʴ�1�u�x�u�?�}����������C�����0�9�;�u�$�5���Y����J��R�����u�=�u�0�8�$�}���Tӑ��[F��RN��4���0�&�;�_�w�.����<����QF������0�;�4�1�$���������lǻC�����
�u�$�4�6�8����Y����[	��h�����4� �u�&�6�<���������X��U���'�!��u�$�/����:����F�A�����&��1�0�$�.�6�������9F��F*�����:�,�o�0�#�)�W���ݣ��R��R������|�u�u�'�/�W���Y���F�d�����>�-�h�u�6�-����J���F���U���
�:�<�_�w�}�W�������F�
P�����4�;�u�u�w�}�ZϷ�Yӕ��l
��^�����'�d�u�:�9�2�G�ԜY���@��^�����h�u�&�'�#��4���U�������*���<�_�u�u�w�.����
���X��D/������y�u�u�z�4�Wϭ�����Z��R����1�"�!�u�~�}�W���
����R)��N��Kʦ��!��!�%�t�W��Y����@��[�����6�:�}�b�3�*����P��ƹK�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���_�u�x�1�#�}��������_F��^ �����=�u��a�]�}�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���lǻC�!���6�;�'�9�;�3�Ͽ�Ӗ��V
��R
����u�:�8�!�?�)�Ϯ�	����VF��[��U���u�3�!�0�6�>��������[��d��6���4�0�:�!�8�.�}�������@N��Z��6���-�_�u�0�>�W�W���Ӕ��Z��R
��]���%�0�9�f�~�)��ԶY���K�`��ʐ�4�9�_�u�w�}��������G*��R�����!���n�]�}�W���Tӧ��A��=N��U���&�1�'�&��)����Dӕ��W��D��N�ߊu�u�u�x��)�W������F�C��ʡ�<�u�&�!�2�;����4����]F��RN�����u�0�4�u�6�<����Y����]F��C��U���u�x�u�u�.�1�Ϫ�Y����V��C�����=�u�<�0�>�8���� Ӊ��G��r�����8�'�_�u�w�}�Zύ�5����[��^��ʻ�0�0�u�;�#�8����Y����[��v-��U���4�&�u�=�w�<����Y���F��X�����u�=�u�=�>�}�������F�N�U���:�=�#�u�>�8����Y����V��QN�����4�<�u�:�:�)�Ϫ�Ӣ��^��d��U���x�u�;�0�9�1�1���s���F�������;�=�<�u�?�3�W���Y����@"��V8�����,�i�u�&�6�<����=�����Y��E���u�&�4�4�6�4�>��Y�����Rd��U���u�&��!��1����Y����@"��V8�����,�c�1�"�#�}�^���
����R0��^
��U���e�e�n�u�w�}������ƹF�N�����<�n�u�0�3�-����
ӥ��P��t�����n�_�u�x��.�W����ƣ�G��DN��U���u�0�!���4�W���Y����]l�D������!�u�u�k�}��������G*��d�����1�0�&� �w�}�K���
����V��B���ߊu�&�4�4�"�}�W���Y����@"��V!��&���_�u�&�4�6�<���������V������,�f�n�w�.�6�������W)��R�����!��9�1�;�u�^�Զs���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�u�:�3�>�4����8���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���_�u�0��3�8��ԜY����V��d�����>�-�_�u�2�4�}���Y����Z��P1�����4�%�0�9�d�t����s���F�������;��0�&�p�z����s���F�D�����'�i�u�&�8�;����s���F��DךU���u�u�&�4��9�W��
����\��h�����&��1�0�$�3�L���Y����]��QUךU���;�u�3�_�w�3�W�������`��S
����_�u�x��2�8�����Ʃ�G��T��ʺ�u�0�4�u�9�.�%������P	��V��U���u�x�u�&�3�/��������F��
�����,�3�'�!�2��3���4����JO�@��ʢ�9�u�4�0�w�p�W���Y����U��R ��U���:�0�6�6�2�?����Y����W��N�����<�u�6�:�9�8�W���s�����V �����u��:�u�?�}����	����Z��S������a��u�;�>�Y���s���E��\1��0���0��8�'�]�}��������A�������"�'�{�$�8�;���� �Ξ�OǻN�����8�%�}�u�w�}�$������� �	N������>�-�u�z�}��������T��N��Uʦ��0��!�w�`�W�������G�N�U���u�!�
�:�>���������W	��C��\���u�u�&��2�
�W���D�ƿ�p	��`�U���x�u�;�u�#�����s���F��e�����u�h�u�&�6����Y�������*���<�
�0�!�%�l��������9F�N�����3�:�&�u�i�.�4���-����]�N��ʦ�1�9�2�6�!�>����Nӂ��]��GװU���u�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�}�Z���*����F�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�_�u�x�?�2�(�������l�C�����4��>��:�1�4��������X��U���&��!��#�/�}���T����X9��T+��Dʦ��!��9�3�1�_���Y����[	��h��0���u�&�4�4�6�4�3���M���K��X��ʶ�u�&�:�3�8�.�}���T����X9��T>��ʦ��6�8�;�w�p��������v��D�����9�1�9�}�~�}�Z¨�������x�����6�8� �_�w�p����&�Ư�	��Yd��Xǣ�:�>�4�6�9�}��������W"��X��U���#�:�>�4�4�>�������Aǻ+����-�u�;�<�.�*��������F��c"��U���2�;�'�6�:�-�_���Y����u��C'�����u�k�>�<�$��4������F��N�����;�o�u�4�$�W�W�������R�=N��U���9�u�u�u�w�}�Iύ�����_��N��U���u�x�<�u�$�9�������F��vN��U���u�u�k�&��)�8������F�C����&�1�9�2�4�+����Q����\��XN����u�u���w�}�W���Gӕ��R��V��1���f�y�u�x�>�}��������9F�N��0���u�u�u�u�i�.�3���/����w
��G�U���<�u�&�1�;�:����Y����qF�N��U���k�&��0������Y���K�^ �����9�2�6�#�4�2�_������\F��=N��U�����u�u�w�}�Iϭ�=����R
��s��@���u�x�<�u�$�9�������F��gN��U���u�u�k�:�2�q�W���Y���F�C����&�1�9�2�4�+����Q����\��XN����u�u���w�}�W���Gӕ��R��V��1���c�y�u�x�>�}��������9F�N��%���u�u�u�u�i�.�6������F�N��U���<�u�&�1�;�:��������Q��X����_�u�u�u������Y�����T��:���u�u�u�u�w�p����
����\��h�����a�u�:�;�8�m�}���Y�Ư�P��B����u�e�|�u�w�}�W���Y���K��YN�����:�<�_�0�3��;��