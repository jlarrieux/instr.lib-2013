-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����E��[�����,�6�:�;�2�s��ԑTӧ��[	��*��U���0�u�;�u�8�8�4�����ƴF��^	�����'�?�6�o���(��L���"��RT��Dʔ�2�&�u�e�e�p�}��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�d�U¶�u�e�g��'�/����7����]��~ �����;�&��'�8�<����T�ƍ�_F��P��U���0�#�1�x�w�<����ӯ��G��R ��U���0�;�9��1�/�������K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X�߇x�x�u� �'�.�Mϊ��Ư�^��R �����0�0�!�u�w�2����Y����
��DN�� ʦ�;�=�:�<�2�p�W���Y�����VN��U���4�!�'�6�8�6� ���Ӏ��B��T��ʴ�8�9�<�9�w�;����T���F�N�����&�:�<�<�6�}����W���F�N��U���u��0�6�8�6����Ӓ��@��^�����3�0� �;�.�/��������Cl�N��U���u�7�!�0�9�����Ӈ��)��E-��[���_�x�u�u�w�}�W�������B��DN����=�u�<�<�0�8����Ӥ��V%����U���'�8�;�&�5�}�}��Y���F�R��ʚ�0��>�6�4�8�W���Y����VF��C�����;�u�0�6�2�W�Z���Y���F��A������6�:�u�w�q�ϰ�Ӕ��Z��R
��U����&��>� �1�W���	����K�N��U���!�0�0�:�2�2����Y����@F��T����u��0�!�:�3�W�������Q��@GחX���u�u�u�u�w�2����Y����@F��Z�����&�4�!�'�6�8����ӄ��@��R
�����6�9�{��%�3�}��Y���F�C��ʡ�4�&�!�:�w�$��������G0��^
��ʳ�9�0�u��"�)����ӄ��\��=C�U���u�u�u�'�2�*����:������D�����;�u�!�'�$�>������ƴl�N��U���u�:�4�0�;������ƥ���RN��ʶ�6�0�7�3�%�}����������RN��U���0�9�{�x�w�}�W���YӉ��@��\+�����!�6�;�7�w�.�Ͽ�Y����]��RN�����u�:�u�;�w�/����s���F�N�����u�0�1�u�8�/�����Ǝ�@��\N�����&�<�u�=�w�+����Y����Z��^	�����u�u�u�u�w�8��������V��u��6���'�&�;�u�3�8�}��T���F�N�����:�9�"�;�w�4����Y����@��C�����&�2�4�&�1�/�ϵ�����\��Y	�����'�x�u�u�w�}�Wϱ�Y��ƴF�N��U���u�u�u�u�w�}�W���&����l9�N��U���
�
�
�
�w�}�W���Yӹ��l9��hd�U���u�u�u��$�����Y�Ɠ�OF�N��U���
�
�
�)�w�}�W���&����l9��N��U���)�
�
�
��W�Z���Y���F�N��U���u�u�u�
�w�}�(���Yӹ��F��hN��U���u�u�
�u�w��W���&���l9ǶN��U���u�u�#�'�;�}�W���&���O9��N��*���)�
�u�)��}����YӚ��OF��h1��U���)�u�
�_�z�p�W���Y���	��B ��U���u�u�)�u�w�!�W��������N��U��u�u�g�u�w�m�W���H�ư�T�Kd�U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u���(���&����l9��h1��*���
�
�
�
��W�Z���Y���F��X��#���1�u�
�
���(���&����l9��C��U���u�u�u�u�w�}�W���Y���F�N��U���
�
�u�u�w�}�W���Y����lF�N��U���u�
�
�
�z�}�W���;����_��P�����
�
�
�
���(���Y����l9��h1��*���u�u�u�
���(���&���F��C��U����!�o�:�6�8��������GF�� ��U���'�;�0�1�w�2����Ӏ���������<�0�7�3�%�W�Z���Y���F�X-�����9�1�4�&�%�.�W���Y����C
��^��:���6�:�>�;��>����Y�Ƹ�VF��E��X���u�u�u�u�w�2��������V(��CN�����4�%�;�4�#�/��������Z��D�����_�x�x�u�w�}�W���-����F��C�����f�'�&�;�w�9����Ӥ��V%�������0�6�:�<�>����s���F�N�����'�'�&�!�3�<����
Ӓ��@�������,�_�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��s���Q��NN����u� �0�<�2�s��������W����N��� �0�<�0�y�(����&����R
��=�����u�:�>�_�w�.�W���ݶ��w��V�����&�u�:�>��:��������@"����N���;�<�,��2�>��������P%��Y��U���2�;�'�6�]�}�8�������u��X��U��<�u�;�0�2�}�J��s�Ƨ�\��z�����!�u�u�o�>�}�������U��U�����_�u��&�#�}�W���Y���F�N��U���9�4�n�u��.�4���Y���F�N��U���;�&�1�9�0�>�}�������XF�N��U���u�u�o�<�w�)�(�����ƹ	��B ��U���u�u�u�u�w�}�W���Y����T����G���&�}��0�4�2�������W	��C��\�ߊu�� �!�6�4�W���Y���F��X�����0�;�_�u��.�4�������K�N��Oʺ�!�7�:�0�9�f����6����_	��^ �����:�;�0�n�]�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���l�:��U���4�0�,�<�w�4����s���W�c�����u��0�0�.�>�����Ƹ�VF��D��ʱ�8�<�{�x�w�}�^Ϛ�����G��R
��ʺ�u�=�u�:�0�4�Ϙ�W���F��*�����=�u�1�0�3�)����Ӗ��@��Y��ʶ�6�0�u�:�'�2����Y����Z��[�����u�u�u�=�w�2����UӇ��V��X-�����9�1�4�1�w�(����;����_��P�����x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z������P��RN��9ʺ�u�#�'�9�4�4��������G��^ךU���;�9�7�:�0�8����Y�Ʈ�\
��YN�U���&�n�u�x�w�8�����Ƹ�VF��M��ʡ�0��u�=�>�s�W��Y����R��C�����u�:�<�u�>�5�����ƪ�\��_�����9�6�u�:�6�3�Yϝ�����X��N�U���0�u�<�<�0�5����Ӌ��GH��_�����u�0�;�0�w�)����Ӓ�� �������6�_�u�x�6�}�����Ƹ�VF��P	������_�u�<�9�1��������F�T�����4�u�h�3�;�8�}�������	��P	��3���%�u�u�:�;�<�W������l�C�����0�4��<�#������Ƹ���R��ʱ�9�,�1�#�%�4����Ӓ����RN�����<�;�_�u�z�u�Ϻ�������[��ʡ�:�3�<�u�;�-�W�������	�������1�u�;�0�>�:�����Ɵ�Z ��N�U���<�!�'�4�$�:����P����\��V ��U���9�,�=�<��'�W�������AF��"�����}�y��0�4�2�������9F��^	�����u��2��#�>�'���Y�Ǝ�\
��Y8�����>�0�4��6�3����T���W	��C��\���u�u�u�u�w�}�W���Y���F�T��]���0�&�k�3�;�8�L���T�ƣ�W��R�����0�e�u�<�;�-��������J�������u�<�<�2�2�:�W���;����_�N�U���&��>�1�2�8�ϭ�����C��RN�����9�6��6�8�}�W��� ����
��R����0�:�0�"�]�}�Zϰ��Ƹ���A��ʳ�:�u��2��)����	�Χ�E��[��3���:�u�u�|�w�5�W���Y����R��Yd��X���&� �0�u�8�5����Y����@F��R�����'�9�6��4�2�W�������G��]�Uʶ�;�!�;�u�<�<����<����V��Y
��U���;�0�0�_�w�}�W���Y���F�N��U���u�u�u�u�m�}��������X ��C��X��u�:�u��2�>��������l�C��6���!�<�u�0�#�/�����Ư�\��T��ʴ�!�'�:�4�2�1�2���7����C��R�Uʶ�;�!�;�u�<�8����:����z��ON��U���;�0�0�_�w�}�W���Y���F�N��U���u�u�u�u�m�}��������X ��C��X��u�:�u��2�>��������lǻC�6���!�u�:�4�w�4����Y����\��B�����<�9�'�4�w�3��������^	��[�Uʦ�2�4�u�u�8�2�������F������1�:�:�;�p�<����C����G��DN��U��|�_�u�<�9�1�W���:����e��S"��U��7�:�0�;�m�}����B���K��E��ʦ�;�u�0�0�w�4����W����Z��[N��U���4�9�
�&�w�}�W������R�
N�� ��u�&�2�4�w�}�������F�N��Oʷ�:�0�;�o�w�/��ԶY���g��x�����>�;��;��(��������VF��R
��ʸ�;�u�:�%�9�3�Ͽ�Y����@�������x�u�=�'�9�}��������_	����U���0�u�;� �$�}��������V��_�����9�u�:�9�w�<�}���TӋ��T��[�����#�'�9�6�>�:��������AF��C��U���2�0�6�8�8�8�Ͽ�Ӓ����N�U���;�6�u�!�w�(����Y����u��YN�����<�!�;�u�;�>�ϱ�Y����u6��N��U���<�_�u�x�#�4�W���������GN����� �0�u�=�$�*��������F��R��ʡ�8�u�=�_�w�p�8�������Z��N �����0�u�&�<�$�<�����ƭ�]��X-�����9�<�u�'�6�8�Y�������Q������&�'�;�n�w�<��������V��X��6���!�6�o�&�0�<�W���[����]ǑN�U���0�6�8�:�2�)�W���Y����]��XN�����8�9�<�9�w�4����WӢ��E����U���,�&�2�4�$�}�Z�������C
��^ �����'� �<�2�:�/�W�������GHǻC�!���8�-�3�;�"�}��������R
��@N�����;�!�;�0�8�}��������]��Y�� ���'�!�_�u�z�>����Y�ơ�K��ZN��ʺ�!�3�'�:�8�3�Y�������Q����*���:�!�u�!�>�:�}�������F��Z����� �u�3�:�8�3�;���Cӕ��]��^��6���!�4��;�"�f�}������K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�u�x�u�~�����Y�Ƹ�T��(��Uʁ�<�u�&� �2�}�ϭ��ƻ�V��u��6���0�2�u�&�>�}��ԜY���F��R��ʱ�8�<�_�u�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���F��P	��3��u�%�:�0�$�<����UӤ��V%��N�����0�<�_�u�w�;�����Ƹ�VǻN��U���4�9�u�u�k�}����B���F��r �����&�i�u�4�$�f�W���Yӄ��T��q��I���4�&�n�u�w�8��������T9��P�����9�|�!�0�]�}�W���<����V9��R�����n�u�u�u�5�3����Y�����V��*���_�u�u�u�z�
�W���^�ƻ�]��c�����u�:�6�4�0�}��������JF��CN��U���&�!�!�u�!�4�}���Y�����V�����!�u�'�7�2�.�}���Y�ƥ���V��U���;�u�u�u�w�?�������F��CN�����0�3�_�u�w�}�������F��SN��N���0�1�%�:�2�.�#�������9l�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�u�z�}�^Ϛ�����G��R
��ʺ�u�=�u�:�0�4�Ϙ�W���F��*�����=�u�1�0�3�)����Ӗ��@��Y��ʶ�6�0�u�:�'�2����Y����Z��[�����x�u�u�=�w�2����UӇ��V��X-�����9�1�4�1�w�(����;����_��P�����u�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��Yӥ��]��d�����0�&�4�0�2�q�8���:���Zǻ���ߊu�u�3�4�2�8�W������F��c�����u�u�u�u�j�;����s���F��X	�����<�0�u�i�w�<���Y���	��P������%�}��0�����)����[��
�����d�u�h�}�#�8���Y����VO��N��Uʺ�4�0�9��0�����DӀ��@��N��Uʺ�:�;��9�w�}�W��Q����A�	N��R��u�u�u�:�8�3�!�������[��V��N�ߊu�u�9�<�w�4��������|��t��U���;�u�u�u�z�}����������V�����&�0�u�=�"�9��������WF��X�����,�!�0��;�3�}���Y�����[���� �0�!�0�w�/�W�������P
��\N�����&�_�u�u�w�	����?���F�������n�u�u�w�2��������C�
N�����0�3�_�u�w�}�Z�������VF��^�����&�o�:�1�2�8�������F��������u�:�u��:����)����F�N�U���%�2�!�u�9�8��������V��_�����=�u��2��)����	�Ɗ���^ �U���u�:�1�0�2�8����ۉ��T��C��%���r�<�=�1� �)�W���Y����v��s�����%�}��2��)����	����T�_�����:�e�n�_�w�}�W��:����VF��RN�����9��2��/�s�>�������VF��B�����3�'�:�0�4�>�����Ư�P
��N��U���u�0�:�0�#�8����Y����p
��E�����1�0�_�u�w�}�5���:����T��O��Hʺ�1�0�0�0�#�4�ǵ�����X#��R �����0�|�_�u�w�}�Z��������������{��&�4�#�4�W���IӇ��V�������0�2�u�3��.�4���Y�����X+�����0�!�<�0�<�8����:����z��OG�����u�u�u�u�8�2�������F�F�����u�k�r�r�l�}�W���YӉ��F��V��9���i�u�'�0�]�}�W���T����|3��r<��!��� �t�:�:�9��Ͻ�����@��CN�����4�0�,�4�#�/�������F�C�����0�!�u�0�6�.�W�������V��^�����:�:�;��;�9�����ƪ�_��@�����u�u�x�u��:����Y����Z��[��U���&�u�=�u�$�3��������V�������{�u�u�u�2�.�ϱ�����R
��{�����_�u�u�u�w��������	��B �����u�n�u�u�w�8�Ϸ�B����������;�u�'�6�$�}������ƓF�*�����4�u�1�0�8�}�#�������9F��r
��1���6��%�}�~�a�WǱ�����u ��X��!���9���%�~�W�W��Y����T��_�� ���!�_�u��"�)����Y����p	��C8�����9�_�u��"�)�W���Y����p	��C"��N��1���_