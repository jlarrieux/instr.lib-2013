-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����A��s�����9�6��%��s��ԑTӧ��[	��$��ʔ�8�'�4�_�z������Ɯ�\��CT��-���`�a��x�w�<����HӬ��JF��_חX���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z�������W��X�����u�4�<�;�;���������%��G�����_�x��9��:��������VǶN�����4�u�;�!�"�8��������R
��Y�����:�_�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��s��ƴF��E�����=�&�3�9�w�4��������_��DN�����=�u�!�
�8�4�W����Ƹ�R��_חX���u�u�u�u����������(��RN�����0�u�:�!�2�3�­�����Z��X��U���!�0�x�u�w�}�W���?����w��E������%�_�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���9l��U��ʼ�0�y�"�'�l�}��������@��[����c�{�9�n�w�(�Ϸ��Ȣ�^��T1��Ĵ�9�_�u�&�w�2��������Z
��^�����9�n�u� �2�*����������d�� ���"�'�{�>��<��������Z��X����_�;�<�,��<����)����_	��c��9���&�u�2�;�%�>�}���Y����F��Z������6�0�o�>�}��������W��N�����'�9�6��4�2�W���ӏ��V��T��F��u�%�'�}�w�}����	����@��N��U���
�:�<�n�w�}�$�������\��YN�����2�6�_�u�w�+����Y�ƥ���h����u�u�&�&�%�8����Y����G��X	��N�ߊu�u��4�2�3��������Z��C
�����
�0�!�'�e�}�������F�_����2�'�7�!�]�}�W�������_��^ ��:���o�<�u�!��2��������Q��X����n�u�x�m�o�}�Wϭ�
����p	��QN����!�
�:�<�l�W�W���*����c��R8�����u�;�&�1�;�:��ԜY�ƿ�G��g����<�u�!�
�8�4�(������F��@ ��U���u�x� �f�f�W�W���
����z��[��Oʼ�u�!�
�:�>�f�W���
����z��T��ʦ�1�9�2�6�!�>����Nӂ��]��G�X���d�{�_�u�w�����0����Z��C
�����
�0�!�'�f�}�������K�d_�D���u�&�4�4�9�m�MϷ�Y����_	��T1�����}�b�1�"�#�}�^���Tӵ��WǻN��1�����u�u�9�.��������V��EF�U���;�:�e�n�z�}�F���s���@4��S/�����u�u�;�&�3�1��������AN��S�����|�u�x� �g�l�}���Yӕ��P��B�����o�:�!�&�3�1����s���@'��B�����u� �u�!��2��������R��S�����|�u�x�u�c�s�}���Y����F��C?��U���u�!�
�:�>���������W	��C��\��u�x��`�g�8�Ϙ�����P6��T,�����%��n�_�%�5��������g*��QN�����0��:��8�6����/ӏ��9F�N�����u�;�4�'�.�)�W���ӕ��G��N��ʴ�'�,�&�/�w�.�W��Y����A��R
��ʡ�0�8�-�8�:�3����Y����c%��B�����_�u�x�:�w�5�W���7���@��V��1����'�,�;�w�}�����ލ�A��CF����!�u�|�_�w�4����
����r��N'��U���<�;�1�m�%�<�(���Y����G	�UװU���#�:�>�&�0�)��ԜY����R
��v������<�;�1�w�4����M�ƨ�D��^����<�;�9�&�4�(�8���*����W\��^	����u�:�;�:�g�f�Wϭ�����@'��B�����<��:�o�5�2����s���E��\1�����_�7�2�;�]�}�Zώ��Ƹ�VF��C��U���u�;� �&�>�)�W�������F��[�����<�&�_�u�z�6����*����V��E-�����9�8�;�&�>�}��������D�������0�!�1�u�z�}����������V��ʠ�;�6�&�4�.���ԜY����R'��V��<��u�&�2�0������0�����Y�����4�;�e�|�]�}�3���8����z��S�����0�}��!���^��
����WN��V����|�_�u�x�?�2�(�������V��X�����:�_�u�x�?�2�(���5����R4��R�����:�0�;�4�!�-������ƹK��_��*��� �0��&�#�)�(�������@3��E<�����u�x�#�:�<�<����
����A��Y�����;�1�&�=�$��������F�A�����&�4�6�,�;�.����6����]��Y�����6�,�9�&�>�(�8���s���E��\1������!�:�3�w�2��������f��[�����_�u�x�=�8��W�������R��V��U���7�:�0�;�$�)��������_��=N��X���:�
�u��6�)����Y����T�������=�&�|�u�z�+����ӕ��G��a��ʡ�
�:�9�4������/����l�C�����4�&�4�4�9�}�3���8����z��\'�� ���8�9�&�0��>���Hӂ��]��GךU���=�:�
�u��)�>���
����r��N'��]���%�!�4�%�2��������F��@ ��U���u�x�#�:�<�<��������V��B �����}��4��3�8��ԜY�˺�\	��VN������!�4�<�w���������Z��XךU���=�:�
�u��>����0ӕ��P��B�����1�u�x�#�8�6�ϭ�����F��D/�� ���!��2�0�]�}����=����\��X�����u�;�<�,� �/�Y�������c��u�����u���_�w�}�����ơ�CF�N��Uʾ�;� ��8�;�.�������F��Y��&���9�&�0��4�8�W��Y���Z��P��O���_�u�u�u��8��������\�N��H����0�6�:�<�<����Y���F���U���0�0�u�h�d�}�WϮ��ơ�CF�N��Uʴ�#�%�4�0�2�}�W���Y���G	��X�������2��$�)�[���Y���F�N��U���u�u�u�u�z�4�Wϼ�Y���5��G�����u�u�u�u�w�c�$�������F�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�;�u�_�w�}�W�������F�N��U���h�u�#�'�;�q�W���Y���F�N��U���u�u�u�u�w�}�W���Y���K�^ �����u�u�&�&�%�8����Y���F�	N��*���9�4�}� �2�����U���F�N��U���u�u�u�u�w�}�W������9F�N�� ���9��0�3�w�}�W���GӒ��Q	��R������!�:�3�~�}�W���Y���F�N��U���u�u�x�u�9�}�}���Y�ƿ�[��~ �����!�u�u�h�w�3����ە��R��Y�����|�u�u�u�w�}�W���Y���F�N��Xʼ�u� �u�u�w�.���� ����~��D!��U�� �&�2�0����������Z��x ��Y���u�u�u�u�w�}�W���Y�����ךU���u��4�!�?�.�!������X��X1�����;�&�!�'��<�������F�N��U���u�u�u�u�w�p�W���Y���F�D=�����4�0�u�u�w�}�J�������V��d�����&�|�u�u�w�}�W���Y���F�N��U���u�x�<�u�"�}�W���
����z��[��U���u�u�k�!��2����Q����R/��V��\���u�u�u�u�w�}�W���Y���F�C�����_�u�u�u��)�>���Y���F�N��U���!��'�,�9�u�>�������_��R�����x�d�1�"�#�}�^���T�ƥ�F��N��Uʦ�4�4�;�u�w�}�W���Y���@"��V/������>�;� ��0��������_�_�����:�e�y�u�z�4�Wύ�Y�����V
�����&�u�u�u�w�c��������@4��S/�����|�u�u�u�w�}�W���Y���F�N��U���u�;�u�_�w�}�W�������G0��^
��U���h�u��6�:�(�!�������F�N��U���u�u�u�u�w�}�W���Y���K�X�����u�u�&�6�"�����Y���F�	N������!��2�2�q�W���Y���F�N��U���u�u�u�u�w�}�W������9F�N��4���8� ��u�w�}�W���Gӕ��P��B�����1�n�u�u�w�}�W���Y���F�N��U���u�u�x�u�"�}�}���
����^)��a����u�:��1�8�4�_�������G0��^
�����_�u��6�:�(�>��Y����_	��T1�����}��6�8�"�������ƹ��T�� ���i�u�!�
�8�4�(�������r��Z!��$���;�1�n�0�3��;��