-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����B%��Q#�����#�1�x�u�"�5�����Ǝ�X��C�����;�9��:�2�)�W�������4ǶN����g�u�0�0�5�/�E��s��ƴK�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���_�x�}�|�e�l�W��� ����GF��C�����;�!� �0�#�}��������]l�/��U���=�&��&�%�8�}��7����]��~ �����;�&��!�%�<�W�������Z	��C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�]�p�'�������g�������;�u�8�9�:�3�Ͽ�H�Ʈ�GJ�
�����<�!�<� �2�}��������9K�N�����{�_�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T��Ɠ9
��E��U���0�_�u�&�w�8��������Z��X����_�u�&�u�2�8��������G��[����&�;�=�&�$�)��������U ��^��������_�$�}�9���4ݰ��^��R ��[���n�x�u�,�#�8��������R��X װ���!�u�$�:�1�8�������C	��d��&���9��>�-�w�g��������T��=N�����3�4�4�u�w�}�ϭ�����Z��R����u�:�;�:�g�f�Wϭ�:����VF�N��U���&�1�9�2�4�W�W�������AF�N����!�
�:�<��8����Hӂ��]��G�Uʦ��0���'�}�Mϱ�ӕ��l
��^�����'�d�u�:�9�2�G���B����#��X�����,�_�4�6�>�8����Y����\ ��F-�����:�,�<�_�w�>��������r+��o_��U���2�;�'�6��}�W���0����	F��C1�����}�d�1�"�#�}�^��Y����V��^��N���u�%�'�u�]�}�W���Y�ƣ�GF��S1�����n�u�u�u��}�W���
����_	��TUךU���u�d�o�<�w�)�(�������F�N��U���;�&�1� �8�4�L���Y���� F��^ �����9�2�6�_�w�}�W��Cӏ��@��B����u�u�u��m�4�W���&����Z��N��Uʂ��u�u�;�$�9������ƹF�9��Oʼ�u�!�
�9�0�>�L�������\��Y��N���x�#�:�>�$�:����s���E��\1�����_�u�&�2�6�}��������\��N�����2�6�#�6�8�u�@Ϻ�����O��N�����u�&�4�4�"�����Y����_	��T1�����}�b�1�"�#�}�^��Yۉ��V��	I�\�ߠ7�2�;�_�w�8�%���C����\����Eʡ�u�b�2�;�%�)�}���Y����[	��<��F؍��u�u�x�!�2����0����kD��^�E���u�u�x�#�8�6�ϩ��Ɵ�^��t�����u�x�#�:�<�<�ϭ�:����R��~GךU���x�=�:�
�w�8��������F�C�����4�4�u�&�6�����P���K��_��*���d�&��8�3�/�F�ԜY���E��\1�����e�_�u�u�z�5����Y���AǻN��X���:�
�u�a�p�z�W���Tސ��\�������4� ��8��t�W���+����kW��N��8���d�_�u�u�w�8����Y����l�N��Uʜ��u�k��g�m�G��[���F��N�����6�:�}�d�3�*����P���kD��^�E���u�u�u�%�%�}����s���F�xN��U��&��!��#�2�Ǘ�U���	����*���2�6�u�u�w�}�6���Y����@4��v
��]���u�u�u�x�w�3�W���&����ZǻN��U���d�u�h�u�$�<�6���Q���F�C����&�1� �:�>�W�W���Y�ƍ�F�	N��R���u�u�u�u�w�}�W������G��[�����u�u�u��w�}�I���^���F�N��U���x�u�;�u�#��������F�/�U��u�e�y�u�w�}�W���Y���F��N�����:�<�_�u�w�}�W���Y���@��R�����|�u�u�u�z�4�Wϭ�����T��N��U�����u�k��0�������F�N�U���u�!�
�9�0�>�W���Y����vF�
P�����3�0�n�u�w�}�W��Y���@��B���ߠu�0�1�2�9�/��������@]ǑN�����3�_�u�'�4�.�_���	����XU��=N�����_�u�u�3�%�.��������R��R-��F���!�0�_�u�w�}��������P
�
N��1����!�:�7�]�}�W���Y����F��SN�����&��;�9�1�W�Wϭ�:����\"��R�����!��!�6�l�W����-���