-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����B"��V���߇x��!�:�m��Ϝ���ƴF��^	�����'�?�6�o���(��L���"��RT��Bʟ�;�4�,�g�f�W�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�CחX���|�g�d�u�8�$����Y����\��'�����0�!�u�:�'�/����s����_
��^	��ʇ�&�'�0�_�z������ƅ�@��Z��ʜ�!�'�4�u�9�2�������K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�_�x��>�}��������Z��V �����u�u��a�{�>��������U	��VN��6ʳ�;�!�:�{�w�)��ԑTӄ��[F����U��6�8�4�<�;�s�Z���Y�Ɗ���YN��X���u�u��:�w�W�Z���HӠ��\��d�U���u�0�_�x�w��%���T���cI��X��I����~�6�;� �8�W�������R��^��U���:�0�w�e�g�m�U��Y�Ɯ�c��CN�U���6�;�u�"�2�}�6�������V[�B�����0�w�e�e�f��Z�ԑT���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C���7�4�,�<�2�f�Wϫ�ӏ��VH��S1�����d�c�{�9�l�}��������]��E�����4�9�_�x�w�$�����Ƹ�R��V������7�4�,��1��������l��U��ʀ���n� �2��>���W����C	��Y��4���_�x�&�;�?�.�Ϫ�����G��Ydװ���!�u�$�&�c�}����YӁ��V��d��Uʾ�<�&���6�3�W���Ʈ�\
��YN�U���&�u�n�u�'�/�_���Yӥ��F������9�2�6�_�w�}�6���Y�ƥ���h�����0�!�'�d�w�2����I��ƹF��r ��U���;�&�1�9�0�>�}���Y����F��^ �����:�<�n�u�w�>�W���Cӏ��@��[�����6�:�}�b�3�*����P���F��Y#��Oʼ�u�!�
�:�>�f�W������\��B�����:�<�
�0�#�/�C�������V�=N��U����u�u�;�$�9�������F��T'��Oʼ�u�!�
�:�>���������W	��C��\�ߊu�u���#�g����
����\��h�����a�u�:�;�8�m�L���YӅ��P��[��U���;�&�1�9�0�>�^����Ɖ�w��Uװ���=�!�6� �2��;ϱ�Y����CR��^װUʶ�8�:�0�!�3�-�O�ԜY�ƫ�]��TFךU���u�����}�W���Y�����R	��U��d�_�u�u�w��:���+���F�N��U���0�0�u�h�f�W�W���Y����F�N��U���u�u�u�;�2�8�W��H���F�v;��'���������#���Y���F������u�h����W�W���Y����a#��c1��!���������>���Cӕ��Z��S��8����n�u�u�w��>���-���F�N��Oʦ�'�;�u�h�u��2���B���F��t/��'���u�u�u�u�w�g�������F��=N��U�����u�u�w�}�W���Y����]��R��H��_�u�u�u���"���Y���F�T�����2�o�u����U�ԜY���p'��n'��0���u�u�u�u�w�3����Y���l�N��6��������}�W���Y����T��S��N���u�u���w�}�W���Y���F��^ �����o�u�n�u�w�}�:���Y���F�N��U��7�!�#�6�8�}�Jφ�J����u ��q(��N���u�u���w�}�W���Y���F��^ �����o�u�n�u�w�}�:���:����z(��pN��U��<�!�2�'�m�}�L���Y����c+��r<��U���u�u�u�o�>�)����C����9F�N��4����u�u�u�w�}�W������V��EN�U���e�e�e�e�g�m�L���Y����a#��N��U���u�u�u�o�>�)����C����9F�N��0�����u�u�w�}�W��
����TF��L��&���_�u�u�u���6���+���F�T�����2�o�u����9��Y���5��h<��;������u�m�.����Y���`#��z/��W�ߊu�u�u����2���Y���F������o�u���u�W�W���Y����~3��N��U���u�u�u�!�>�:�M���4����`D��N��Uʀ�������#���Y�ƿ�A��T��W������w�]�}�W���*����~"�N��U���u�u�!�<�0�g�W͑�<���l�N�����u�u�u���}�W���Y���	F��N�����:�<�n�u�w�}�6���Y���F�N����&�1�9�2�4�+����Q����\��XN�N���u�u���w�}�W���Y����Z�D�����6�#�6�:��d��������l�N��4����u�u�u�w�}�W���Y����_	��T1�����}�l�1�"�#�}�^�ԜY���qF�N��U���u�u�u�;�w�)�(�������P��_����!�u�|�_�w�}�W���7���F�N��U���u�!�
�:�>���������W	��C��\�ߊu�u�u���}�W���Y���	����*���<�
�0�!�%�l�W������]ǻN��U���u�u�u�u�w�}�MϷ�Yӕ��l
��^�����'�a�u�:�9�2�G��Y���6�N��U���u�u�o�:�#�.��������V��EF�U���;�:�e�n�w�}�Wώ�0���F�N��Oʼ�u�&�1�9�0�>����������Y��E��u�u�u���	�W���Y���	F��CN�����2�6�#�6�8�u�@Ϻ�����O��N��Uʖ����u�w�}�W����ƿ�W9��X	��N���u�u�����W���Y����\��D�����6�#�6�:��}�������9F�N��4������u�w�g����
����_	��TUךU���u������#���CӉ����h�����_�u�u�u���2���Y���\��YN�����:�<�
�0�#�/�AϺ�����O��N��Uʔ� ���u�w�}�W����ƿ�W9��P�����:�}�u�:�9�2�G��Y���%��e7��&���u�u�o�<�w�.��������V��EF����!�u�|�_�w�}�W���-����z(�N��U���&�1� �:�>�f�W���Yӫ��g5��y!��U���o�:�!�&�3�(����B���F��a+��9���u�u�u�o�8�)��������P]ǻN��U������u�w�}�Mϱ�ӕ��l��P�����u�u�����2���-����F��C
�����6�_�u�u�w��#���=����gF���U���
�9�2�6�]�}�W���<���F�N��U���;�u�!�
�;�:��ԜY���p#��N��U���u�u�u�;�w�)�(�������F�N��4�����u�u�w�}��������\��d��U�����u�u�w�}�W���Y���@��B����u�u�u���}�W���Y���	F��N�����:�<�n�u�w�}�4���Y���F�N����&�1� �:�>�f�W���Yӥ��r4��~ ��U���o�<�u�&�3�(����B���F��r-��9���u�u�u�o�>�}��������P]ǻN��U���u�u�u�u�w�}�MϷ�Yӕ��l��P�����u�u�� ���%���Y����]F��C
�����6�_�u�u�w��W���Y���F���U���
�9�2�6�]�}�W���*���F�N��U���;�u�!�
�;�:��ԜY���a5��{"��'����u�u�;�w�)�(�������F�N��!�����u�u�w�}��������\��d��U�����u�u�w�}�W���Y���@��B����u�u�u���}�W���Y���	F��N�����:�<�n�u�w�}�%���-���F�N����&�1� �:�>�f�W���YӴ��~F�N��U���o�<�u�&�3�(����B���F��d:��U���u�u�u�o�>�}��������PO��N��ʶ�8�:�0�!�]�}�����Ư�V��N����9�2�6�#�4�2�_������\F��d�����4�u���3�}�W���&����P9��T��]���:�;�:�e�l�W����s����r��R�����9�2�6�#�4�2�_�������Z��SF��\��|�n�u�6�'�2���Y����W��N������'�!�;�?�4�W������F�N��U���e�d�e�e�w�5�Ͻ�����_��
I�U���0�w�e�e�g��}�������V9��N�����_�u�0�0�>�}����Y����P��E��H���y�u�u�4�"�2����Y���l�N�����k�g�_�u�w�(��������G��Y1�����u�k�3�9�2�W�W�������@��G�����1�!�6�
�'�4���Yѫ��p.�=N��U���;� �u�k�u��2���U�����D����u�y�u�u�5�8�W���H���F��^ ����u����u�W�W�������]��S�D�ߊu�u�4�'�>�.����Y���l�N�����k�d�_�u�w�<���Y����u ��q(��3���_�u�u�'�0�`�W��Y����F
��V�����2�h�u�y�w�}��������[�BךU���4�!�'�u�i�%�G��I����V��d��Uʥ�0�u�k�d�]�}�W���&����W��h����u������}���Y����^��S�W����y�u�u�$�1�������F��v:��'���_�u�u�&��(���Yѫ��g9��d��Uʠ�0�%�!�0�9�9����Y���})��v:��!���u�u� �0�$�0�W���[����D�G��U���}�u�u�6�<�`�W���U����	N�����_�u�u�u�i�>�[���YӅ�F��C����e�|�_�u�w�<����Y���A�N�����u�k�}�!�2�.�J���I����F�U��U��}�!�0�&�j�}�G���s���C��S����;�_�u�u�6�/�������A��d��Uʸ�9�&�2�<�w�c�P���s���R��CN��U���;�_�u�u�4�(�W�������9F������&�:�!�h�w�-��ԜY�ơ�_��P ����u�%�;�_�w�}�W�����ƹF��V�����0�0�!�h�w�-��ԜY�Ƽ�G��Y
�����h�u�%�;�]�}�W�������[�X��Y���u� �1�'�;�*�J���	����F�T�����u�k�:�0�{�}�WϮ����F��T!��Y���u�:�8�1�w�c��������F�V�����h�u�e�e�u�W�W�������]��S�W��w�_�u�u�2�l�J���<����9F���G��u���y�w�}��������[�_�����u�0�d�h�w�l�[���YӅ��F�I�Y���u�6�6�h�w�l�[���YӅ��R��^ ��K��r�_�u�u�2�}�IϽ���ƹF��R����u�d�y�u�w�>���Y����l�N�����6�'�,�;�j�}�F��Y����@��
P��E���u�u�'�!�;�0����G����l�N�����k�r�r�_�w�}����D���JǻN�����9�4�'�<�w�c�P���s���A��S�R��_�u�u�&�4�/�W���^����F�E��U��r�r�n�u�w�W����-���