-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����A��s�����9�6�{�=�]�p�6�������\��v�����_�x��<�>�<�W�������6��R1�A߇�x�u�4�0�w�l�=���Y����9K��C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�w�>�W��Hӥ��J��_�����;�9��&�%�0����:����A��X חXʔ�9��2�!�w�8�������}��X ��U���!� �0�!�w�3����ӯ��\��C�����x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�Z��Y����\��N�����<�0�6�0�#�.����������T����� �<�&�3�%�)�ϸ�����]��=C�U���u�u�u�1�4�0����Y���9K�N��U���u��<�u�8�(�ϭ�����RF��@N�����4�<�;�0�2�$����Y����A��V�����_�x�u�u�w�}�WϿ�
����F��CN�����=�;�6�9�"�<�Ϫ�Ӏ��G��X�� ����6�8� ���}��Y���F���ʼ�u�4�<�u�?�3��������e��SN�����&�_�x�u�w�}�W���7����R��^�����0�u�;�:�#�8����Ӕ��Z��E��ʴ�&�'�<�2�z�}�W���Y���@"��V'�����u�<�=�#�;�9����Y����w��~ ��$���_�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���Q��NN�����"�'�n�u�"�8����W����_	��T1�C���9�n�u� �2�4��������P9��S@���ߊu�&�u�:�<���������R
��T�����4�9�_�u�$�}����)����f��^�����{�9�n�u�"�8� ���W����A��s�����<�<�;�&�6�1�}���5����A��y'��8�ߊu�&�u�������	����G��[�U���;�<�,��6�)��������P��DNךU���!�_�u�u��.����Ʈ�\
��YUךU��� �0��&�#�}�W�������R��N��&���9��>�o�>�}��������9F�N��U���u�u�_�u�w�����:����\��YN�����;�_�u�u��<��������GF��^ �����;�1�>� ��<����
����\��XN�N���x�g�{�g�w�}��������V��Y�����u�;� �&�0�8�_�������V�N� ���_�u�u�u�$�)��������_��N��U���9�4�n�u�w�.����)����\��YN�����0�}��8�?�.�5���T�ƨ�D��^�U��� �f�d�_�w�}�W���Yӕ��G��a����<�u�:�9�6�f�W���
����z��N��U���;�1�d�u�8�3���B���`W��d��Uʦ�4�4�;�u�w�3����������Y��E��x�u�d�{�]�}�W�������A��~ ��U��� �&�2�0��}�������K�b_�D�ߊu�u�u�u�w�}�W���Y����r��Z!��#���1�o�:�!�5�2����s���@'��B�����u� �u�<�9�9�C�������V�N�U��{�_�u�u��>����(����F��^	����u�:�;�:�g�t�W��Y����l��SN�����0��:��8�6�}������P��RN��9ʺ�u�'�6��4�/�����ƥ�9F�N��U�ߊu�,�0��0�8�Fן� ����@F��E��U��� �4�u�4�0�}�I����ƿ�T��_����!�u�|�_�w�$�ύ�����'��h��ʴ�'�,�u�4�"�<�W������O��QN�����}�b�1�"�#�}�^�ԜY����6��D�����<�u�'�4��3����Ӕ��T�	N�����;�<�;�1�<�(�'�������W��X����n�u�!�%�w�3�����֍�J9��^�����}�;�!�'�;�/����E���\ ��Y�����l�1�"�!�w�t�}��� ����]��Y��G���
�u�&�4�%�$�W�������A��RN�U���3� �&�2�2�u�FϺ�����O��=N�����9�&�=�&��1��������q	��R�����'�>� ��8�8����,������Y��E��u�&�2�4�w���������	F��V�����}��8�'�4�.��������W	��C��\�ߊu�<�;�9�$�>��������A��N�����;�0�!�'�<�(�'�������T3��C�����:�e�n�u�$�:����8����r��N'��U���;�1�m�'��u�9�������@��b ��ʱ�"�!�u�|�]�}����ӕ��P��E��$���2�0�a��$�ǵ�����P��^ �����u�:�;�:�g�f�Wϭ�����@'��B�����4��o��0�8�Cן� ����}��E�����2�;�!�u�8�3���B����Z��[N������!�'�4��g�$�������A�������6�&�<�2�9�)�W������]ǻ�����&�0�1�1�%�.�6��� ����]��Y��E���
�}��8�%�>��������@F��@ ��U���_�u�<�;�;�.��������U/��R�����&��u�u�9�4����K����GN��B�����&�;� �<�$�9� ���Y����F��P ��U���2�0�!�:�1���������@+��T�����;�1�g�'��u�9�������@��b ��ʱ�"�!�u�|�]�}����ӕ��R��S�����<�0�o� �$�:���8����R��X����n�u�&�2�6�}�"�������U ��G��U���9�4��6�8�u�BϺ�����O��NװU���#�:�>�&�0�)��ԜY�˺�\	��D���ߠ7�2�;�u�w�}�}���Tӵ��V��C�����0�!��"�$���������\��^��6ʴ�1��2�0�#�2��������A2��D#��U��� �&�u�x�w�<����ӑ��P��V�����0�u�0�4�2�(����s�Ƽ�\��DF�����y�4�%�0�;�t�Wϼ���ƹF��QF�����|�!�0�_�w�}�W�������\��g��U��}�!�0�&�j�}����P���F�D"�����:�3��1�/�2�#���4���F�
N��*���<�;�1�u��*��������W��X������y�g�n�w�}�Wϭ�����p	��Q'�����'�=�&���t�W������@��R
�����0�!�:�3��9����-����r%��\����u�u��"�$���������\��^��6��u�i�u�:�"�.����QӍ��D��t�����0��'�=�$��E��P���F�D&������0�3�;�2�����
����O�
N��*���<�;�1�>�>�5��������W��X������y�g�n�w�}�Wϭ�����G%��Q�����:��<���l�W������@��R
��=���0�!�:�3��9����-����r%��\����u�u��2�2�)����0����u	��_��4���|�i�u�:�"�.����Q����[��t�����0��'�=�$��E��P���F�=N��U���<�u�<�<�0�8��������p
�������u�x�u�!�>�}��������G	��X������!�:�3�w�.����Y����\	��V �����0�y�"�<�?�*��������VF��N��X��� �0�3�;�8�)�W���Y����\F��CN�����u� �0�9��8�Ϫ�Y����T��R�����;�u�3�<�w�5����s���K��CN�����0�3�9�:�2�}�ϭ�������[�����4�4�0�:�.�/�������g��	�����&�_�u�u�z�5�����ƣ���[�����'�%�2�!�w�5�W�������]F��,��ʓ�9�0�u�:�1�4����
ӓ��WH�N��X���0�!�>�u�3�<����Y����[��D��ʶ�6�0�u�:�'�-����Y����@��T��U���'�1�6�u�?�}�������F������!�;�u�u�?�4�W���?����VF��RN�����:�=�'��w�3����Y����P�������u�=�u��]�}�W��������E��ʱ�&�4�!�7�8�6��������Z ��_�����u�:�u�u�w�}����8����V ��^��I��� �0�9��2�;����
����_��R�����=�2�x�u�8�3���Y�ƿ�@��C-����u�u�u�u�w�}����,����G%��Q�����|�u�=�;�w�}�W���
����@��R������'�=�&��u�^��Y����]��Y�����0�!�:�3��9����-����R��C^�G��u�u�u�0�$�W�W���Y�ƿ�\��C-�����1�-�:��>��4��Y����\9��D������"�&��2�;����?����Z��t^�G��u�u�u�0�3�4�L���Y���F�N��]���0�9��0�1�4���PӒ��]l�N��Uʦ�:�0�!�:�1���������@+��_��I���:� �&�2�2�u�;���
����U ��S�����<��6�9�f�l�^�ԜY���V
��=N��U���u��"�&��8��������g��z/��D���h�!�
�;�>�3�ǵ�����p	��Q'�����'�=�&��f�l�^�ԜY���V��^�U���u�_�u�u�w�;����8����V ��^��L���!�0�_�u�w�}�W�������\��~ ������<���e�}�JϪ�&����T��������0�3�;�2�����
����_��\����u�u�9�0�w�}�W���
����@��R������'�=�&��u�^��Y����]��Y�����0�!�:�3��9����-����r%��\����u�u�;�u�1�W�W���Y���F��QF�����!�:�3��'�u�F�������F�N�����=�&��0�1�3��������~'��G��Hʡ�
�;�<�;�3�6����
����U ��S�����<��6�9�g�l�^�ԜY���V
��=N��U���u��2�0�#�2��������A2��D#��]���i�u�:� �$�:����1����@��R������'�=�&��m�F���s���F��SN��N���u�u�_�u�w�}�ǭ�
����p	��Q>����|�u�=�;�w�}�W���
����V��X��<���-�:��<���F���DӒ��F��P ��]���2�0�!�:�1���������@+��v��Y��n�u�u�u�2�.�}���Y�����P�����3��1�-�8�	����:���[��X1�����0�}��2�2�)����0����u	��_��4��d�|�_�u�w�}�������F�=N��U���3�&�&��#�2����	����O��_��U���u�u�&�<�?�.�4�������K ��c��8���g�u�h�!��3����ۍ��T��C-�����1�-�:��>�����K����l�N�����_�u�u�u�w���������U/��R�����&��}�|�k�}����
����WN��^	�����0�3�;�0��/����8���O��N��Uʰ�1�<�n�u�w�8�Ϸ�B����]��E����_�u�x��'�1����+����W��D��U���0�6�:�>�4�>����Ӆ��C��V�����!�0�!�'�2�>����+����A��[��U���u�;�u�4�4�5��������WF��G�����0�4�&�!�%�(�Ϫ�Ӏ��@��E�����2�7�:�>�w�W�W��?����w��E�����:�!�:�u�$�*����
Ӓ���������<�0�<�0�3�1�ϱ�Y����VF��P ��ʷ�3�'�u�u�z�}��������V��C�����<�&�u�'�4���������A��[��[���%�:�0�&�6�8��������p
��=N�����_�u�u�3�6�8��������F�N�����1�'�&���-�W��Q����A�	N�����&�h�u�e�~�f�W���������^ �����}�4�%�0�;�t����s���F��R�����&���%�w�`��������V��Y>��¦�0�1�1�'�$��'���^����W��X����u�u��4��9�������F��SN��N���0�1�%�:�2�.�}���Yӕ��R��V��4���,�e�u�i�w���������R
��d�����&��'�,�g�}�W���Y����`��C>����u�&�0�1�3�/�������F������1�0�&�;�>�8��������V��Y>��ͽ�2�|�_�u��>�������F�N��H���!�0�&�h�w�m�^�ԜY����F��E��]���u�u�u�h��)����D���O��NךU����0�!�u�?�}����
������CךU���0�4�0�'�4�3���YӀ����YN�����8�'�6�$�4�����ƫ�]��CךU���x�=�:�
�w�/��������f��=N��U���=�:�
�u��/��������Z[��N��Xǣ�:�>�2�>�8�;�:�������P��_ךU���x�=�:�
�w�� ���:����z��O(��!�����&�:�2�)����0����u	��_��4���x�|�u�u�z�+����ӕ��T��C-�����1�-�:��>��4ϭ�����G%��Q�����:��<���4�F�ԜY���E��\1������!�:�3�w�����:����c����U���x�#�:�>�6�.����)����e��SN������9�1�'�6�u�Z���Y�����X��U���4�!�=�&�w���������ZK��=N��U���=�:�
�u��%�:�������F��[�����&��9�1�%�<�_���Y�����X��U���-��6�=�$��ϭ�����A����U���x�#�:�>�6�.��������WF��V�����<�_�u�u�z�5����Y����R/��������u�u�x�!�2����
����z��D*�����_�u�u�x�?�2�(���+����W��D��U���4��1�0�$�/����T��ƹF������u��4��3�8����Y����W'��E��4���,�<�_�u�w�p����&�ƿ�P��~ ����� ��'�,��p�^���Y����[	��h��4���8�;�u��4�0����(ۏ�l�N����>�4�&�6�"������ƿ�P��a�����4�}�|�u�w�p��������r��Z!��9���u��6�8�%�<�>Ƿ�s���K��X��ʦ�6� ��!�4���������R��^GךU���x�=�:�
�w���������r��Z!��4���,�}�|�u�w�p��������r��Z!��$ʦ�6� ��!�%�<�&Ƿ�s���u��C*��%��� �<�-�u�9�4�ϩ��Ȋ�R��R�����<�u���]�}�W�������PF��GN��U���u�u�>�<�$��4������[�^S�U���u�;�u�:�;�<�}���Y���X%��Q�����!�;�0�h�w�p�^���Tӏ����R	�����u�u�:�!�:�-�_���Y�����D��U���u�u�u�u�w�}�W���Y���R4��R�U���u�u�u�u�w�}�W���Y���F�N��Uʷ�:�0�_�u�w�}�W�������V�N��U���u�u�u�u�w�c��������GJ�N��U���u�u�u�u�w�}�W���Tӏ����[��U���u�u��8�;�����Y���F�N��U���h�u�4�%�2�1�[���Y���F�N��U���u�u�u�x�w�3�W���&��ƹF�N��%���0�;�'�8�9�}�W���Y���F�	N������6�0�0�#�}�W���Y���F�N��U���<�u� �&�0�W�W���Y�ƿ�\��C-�����1�-�:��>��4���Gӕ��D��t�����0��'�=�$��_��P���K��YN�����;�u�u�u�w�.����
����U ��S�����<���h�w���������U/��R�����&��}�x�~�}�Z����ƹ�@��=N��U���u��9��4�8�:���
����F�N��U��&�4�6�,�;�.����6���F�N��U���u�u�x�<�w�(����s���F�D;��4���:�3�u�u�w�}�W���Y���X��b�����0�3�<�0�>�q�W���Y���F�N�U���u�:�9�4�w�}�W���
����G6��D�����u�u�u�u�w�}�J���)����e��S/�����x�|�u�u�w�}�W���Y���Z�U���ߊu�u�u�u��<����
���F�N��U���u�u�k�&�?�.�6��� ۏ�J�N��U���u�u�u�u�w�p��������]l�N��Uʦ�0�!�4��6�8�������F�N��U���4�0�4�<��/�Ƿ�U���F�N��U���x�u� �u�8�1����Y�����O�����&��!�u�w�}�W���Y���@6��D�����<�y�u�u�w�}�W���Y���F�N��ʠ�&�2�_�u�w�}�W�������R
��N��U���u�u�u�u�w�c��������_��N��U���u�u�u�u�w�}�W���Tӏ����[��U���u�u�&�4�6�3�W���Y���F�N��U���h�u��!���W���Y���F�N��U���u�u�u�x�w�3�W�����ƹF�N��1�����u�u�w�}�W���Y���F�	N�����;�y�u�u�w�}�W���Y���F�N��U���<�u�&�2�2�W�W���Y�ƿ�V��S
�����u�u�u�u�w�}�W���Gӕ��R��S�����4�}�x�|�w�}�W���Y���K��YN�����;�u�u�u�w�.��������@)��N��U���u�u�u�h�w���������r��NF��Y���u�u�u�u�w�}�Z����ƹ�@��=N��U���u��6�8�9�}�W���Y���F�N��U��&�6� ��%�$�_��P���F�N��U���u�u�x�<�w�.����s���F�D/�� ����u�u�u�w�}�W���Y���X��v�����4��<�d�{�}�W���Y���F�N�U���u�<�;�1�w�}�W���
����^)��a�����u�u�u�u�w�}�J���8����e��S/�����|�u�u�u�w�}�W���Y���\��U���ߊu�u�u�u��>����5����F�N��U���u�u�k�&�4�(�6��� �Υ�F�N��U���u�u�u�u�w�p����
����Wl�N��Uʦ�6� ��!�4��W���Y���F�N��U���6�8�'�4��4�[���Y���F�N��U���x�u� �u�>�3����Y�����T�� ���u�u�u�u�w�}�W���Y���@'��B�����4��<�y�w�}�W���Y���F�N��ʦ�2�0�_�u�w�}�W�������G7�N��U���u�u�u�u�w�c��������r��N?��\��u�u�u�u�w�}�W���TӉ����Y�����;�u�0�0�6�8�0�������A	��Y��N���u�_�u�x��1�����ƪ�]��V�����!�'�:�!�"�.�}���TӨ��Z��C��U���:�9�u�&�w�5�W���������DN��ʺ�u�=�u�6�"�(����W�Ƙ�Z��DN�����0�4�&�_�w�p��������F��R�����;�"�u� �'�/�W���Y����V��Y	�����u�&�d�-�w���������R��N�U���!�'�u�'�w�8����Ӏ����R�����;�:�u�e�/�}����������VN�����8�1�6�8�#�2�W���s����������<�;�&�0�"�1����I����[�\��[���=�u� �u�1�)�Ͽ�
����VF��[�����=�u�u�x�w�<�Ͻ�����Z��DN��U��� �1�d�m�w�	��������G����U���2�&�u�4�"�}�Ͻ�����E��R���ߊu�x�:�!�8�}��������_��EN��U���z�{�`�h�g�o�A���0�ƻ���Y
����� �u�:�!�2�3��������\ �NךU���"�u�0�u�x�m�Bϳ�����\J��RN��ʦ�3�u�=�:�>�:����Y����V��VN�� ���<�&�:�u�?�}��������Al�C�����!�;�u�<�?�<�$��IӔ��A��Y�����_�u��6�:�(�!������@'��B�����'�4�}��:�/��������Z��d����� ��!�u�j�.����6����A�������6�&�<�2�9�)�^��Y����G	�UךU���6�8� ��k�}�6�������A��fF�� ���:�0�&�;��4����Mӂ��]��G�U���u�_�;�u��f�