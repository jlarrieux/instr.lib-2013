-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����A��~ �����0�3�4�6�!�9�Z�������	F��_ �����8�;�x�u�%�:����)����P��g6��*��`�_�x��#�g�E�������V��=C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Wǽ�Y����%��N�����4�<�;�9��.��������\��E���߇x��9��0�)�W�������9K�y�����u�;�!� �2�)�W�������/��X�����_�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z�ԑT���c��X��Uʁ�<�u�<�0�4�1�����Ƹ�VF��Y��U���0�%�9�!�3�>��������@l�N��U���u�u�:�u�6�5�:���s��ƴF�N��U���>�4��&�6�>�W�������V��_��U���3�<�<�;�$�<�ϫ��Ʈ���Dd�U���u�u�u�u�9�)����YӰ��Z��V��ʧ�;�0�3�:�w�}�ϵ�����P��^ �����u�d�_�x�z�}�W���Y���g���� ���"�9�u�4�4�1��������P	��Q�����u�#�'�u�>�8�Z���Y���F�D<������9�u�&�2�)�Y����ƪ�A��T�����0�!�"�9�w�-����T���F�N�����!�6�:�>�4�>��������@4��C��6���u�&�0�!�y�}������ƴF�N��U���>�#�'�9�4�����Y����P	��Q�����u�<�9�4�'�<�W�������V��T�����u�u�u�u�w�}����
����\��D>�����u�&�;�!�%�:�����ƻ�G��e�����9�6�_�x�w�}�W���Yӭ��CF��_��<���;�=�;�0�w�3����+����A��[�����!�u�2�<�l�p�W���Y���F��EN�����0�<�u��2�>����������B�����=� �1�>�2�}�'�����ƴF�N��U���6�;�!�;�w�2�W����Ư�P
��GחX���u�u�u�u�w�}����4����Z
��V��ʰ�0�,�6�6�2�2�ϱ�Y����C	��G��ʳ�9�0�_�x�w�}�W���YӅ��U ��^���߇x�x�u�u�w�}�W���Ӆ��\��C�����!�6�0�3�4�8�ϻ��Ɓ�pF��DN��ʼ�3�'�0�u�a�?�%���s���F�N��U���&�8�8�'�w�)����Q����A��T�����u�u�|��<�<��������G��q���߇x�u�u�u�w�}��������[	����U���u�=�u�:�1�4����
Ӓ��GF��YN��U���9�0�u�,�8�8�Z���Y���F�D������y�!�0�%�.�W�������\��^�����4�0�4�%�>�9�������F�N��U���0�!�:�u�?�}�6�������V��YN�����>�_�x�x�w�}�W���Y�Ƃ�G�������&�4�>�4�2�4��������u��X�����4�u�0�"�2�}��ԑT���F�N�����<�<�;�&�$�2����Ӄ��[F��^	�������u�=�$�2����	ӏ��]��R
חX���u�u�u�u�#�}�����Ƹ�VF��[����� �0�u�!�>�}��������G�������u�=�!�x�w�}�W���Y�Ƹ�VF��E�����3�6�0�!�#�<�W���
Ӊ��	��C��U���%�;�;�u�$�)���Y���F�N�����6�0�!�!�6�}����ӄ��^��^�����<�=�!�0�8�9�������z��C�����u�u�u�u�w�*��������Z�������<�;�u� �w�.��������Z��C�����0�!�4�1�2�.�Z���Y���F�^ �����0�:�,�}�>�5����Ӓ����R�����4�!�'�6�2�;�����ƿ�_��R
חX���u�u�u�u�5�}�'������9K��C��U���u�u�u�=�w�4��������P��CN�����4�0�u�&�6�9����ӄ��G��R�����u�u�u�u�w�}�����Ʈ�G��QN������{�u�=�w�l��������Z��Y��ʧ�4�u� �_�z�}�W���Y����UF��Z��U���"�9�u�&�#�8�F����ƨ�_��C�����0�!�6�0�1�>����s���F�N��U���u�d�3�4�#�2��������UF��_��<���'�u� �!�'�4�ϼ�Y����S��^חX���u�u�u�u�3�1�Ͽ�Ӓ��]F��S�����=�u�'�2�9�1��������]��XN�����4�0�x�u�w�}�W���Y����_��V�����%�9�!�1�4�8�������KǶN��U���u�u��0�$�>��������P��CN�����4�0�u�&�>�8����Ӓ��G��Q��ʰ�6�%�_�x�w�}�W���YӒ��GF��RN�����&� �0�u�8�1����	Ӓ����Q�����u�;�u�0�#�}���Y���F�N�����0�!�1�7�w�m�Wǻ�����\F��RN�����<�!�'�<�#�/��������R
��@חX���u�u�u�u��8����Ӆ��U ��^��U���6�9�!�:�w�8��������[��S
�����,�4�_�x�w�}�W���YӇ��Z��Y��D��_�x�x�u�w�}�W���Y����^��^��U���u�1�u�&�3�4�W���Y����R��Y�����!�:�u�'�w�2�Ϸ�s���F�N��U���u��a��4�0��������[��T�����!�<�u�;�2�/��ԑT���F�N��Uʁ�0�%�%�9�9�}����Y����F��C��U��� �0�<�u�w�$����s��ƴK�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���_�9�7�4�.�4�������9F��D�����&�1�9�2�4�l�A�����ƹ����Ļ�8�'�6�&�3�<��ԜY����D	��>��1���4�9�_�u�$�}����)����R��Y��Ĵ�9�_�u�&�w�2��������G/��R�����<�<�;�&�6�1�}������u��C'�����:�3��9�w�.�WϹ�����l�N�����9�6��6�8�}�W�������V�
N����u��6�;�#�3�������V�=N�����_�u�u��$�)�MϷ�Y����V��=N��U���%�0�9�u�w�3��������l�N�����'��9�u�w�3��������F�D>�����u�u�;� �$�:����Aӂ��]��G�U��� �l�m�u�w�.����6���	�������g�u�:�;�8�m�^���T�Ɵ�H��R ��3���!�;�0�%�8�;�4���B���P��R������u�3��6�)����	����U%��TN�����x�u�4�<�w�+�����Ɗ�P��DN��ʡ�<�u�:� �2�<���J�Ƙ�Z��X
��ʦ�:�9�_�u�z�.��������F��_�����u�4�u�:�w�8�Ϫ�
����/��N��U���6�&�=�#�w�}��������F������;�=�%�!�>�}����������Y	��U���&�%�:�!�>�s�W�������VF��t�����'�4�2�
�w�.��������R��]�����:�g�_�u�z�����Y����A��T�����u�&�<�u�6�:�W�������Q��A-��3���:��;�0�#�W�W��-����R��^�����u�;�,�&�'�2��������R��d�����!�;�u��%�;�8�������\�!�����6�:��;�2�)�W���Y���F�N��U���u�u�u�u�w�`��������X ��C�����x��'�3�w�5�W���������V�����;�!�0��0�/��������^��_�����1�9�,�u�z�}�Ϫ��ƪ�_�c��U��� �0�u�!�2�}����Y�����������,�:�=�'�w�p�W���Ӗ��[��XN�����'�%�'�6�2�;����Ӈ����VN�����0�!�_�u�$�?����:����p��g��1���,�4�2�
�w�.��������R��V�����:�m�_�u�z�����Y����U ��[�����9�,�<�u�9�/��������V��NN�����4�6�<�0�2�<�%������F�:��ʴ�6�<�0�!�%�}����
����A��D��U���2�{�u�6�9�)����/����J%��Q�����%��9�o��8��������w��N<�����_�u�u�u�w�}�W���Y���F�N��U���u�u�h�>�8�;�4���)����V
��dךU���;�9�>�:�1�����Y�Ɵ�EU��E��]��f�1�"�!�w�t�W���Y���F�N��U���u�h��9��8��������JN��V�����6�y�>�#�%�1��������lǻ�����&�0�!�'��1�'���Y�Ʈ�\
��YN�U���&�n�u�&�0�<�W�������A��T�����;�1�}�u�8�3���C����G��DN��U��|�u�x�u�f�s�G�ԜY����R
��e��1����!�o�&�3�1��������AN��
�����e�u�h�}�#�8���Y���l�D������4��!��)����Cӕ��l
��^�����'�f�u�:�9�2�G���D�Σ�[��S�R��n�u�&�2�6�}�4�������]������g�u�:�;�8�m�W��Q����A�	N��R��x�u�g�{�]�}����ӕ��V ��R��U���<�;�1�d�w�2����I����N��_��U��r�r�n�x�w�l�Y��s�ƿ�T�������=�&���'�m�Mϭ�����W��X����u�h�}�!�2�.�J���I����K��\����<�;�9�&�%�>�'�������C��N�����}�d�1�"�#�}�^��Yۉ��V��
P��E���u�x��g�f�}�����ƿ�A��g�����<�0�u�u�>�3���Y����G	�N�Uº�=�'�u�k�p�z�L��Y����l�D������4�!�=�$��'���J����Z��SF�U���;�:�e�u�j�u����
���V�N�U��{�_�u�<�9�1��������@��g��A��&�2�0�}�f�9� ���Y���F��C����u�e�|�u�z��E��s�ƿ�T�������0�!��%�g�g����������Y��E���h�}�!�0�$�`�W��P���5��C�Uʦ�2�4�u��2�;����)����\��^	����u�:�;�:�g�}�J�������[�^��N���u�d�{�`�]�}����ӕ��V ��T�����0�u�u�<�9�9�E�������V�S�����'�u�k�r�p�f�Z���K����F��P ��U���0�3�6�0�#�4����Y����V�N�����u�|�o�u�8�5����G����]�N��D��u�&�2�4�w���������c��N����0�}�e�1� �)�W���C����G��DN��U��|�u�x��f�l�}���������[��U���;�1�f�u�8�3���Y���\��E��K��r�n�u�x��j�Z�ԜY����R
��v
��Oʦ�2�0�}�d�3�*����P���	��R��H���e�|�u�x��o�F���
����_F��X��:���6�u�u�<�9�9�E�������V�S�����'�u�k�r�p�f�Z���K����9F�N�����u�=�!�!�2�-�����ƿ�R�������=�u��u�;�>�W���Y����A��E���ߊu�x�:�!�:�'�Ϸ��Ɵ�U��=N�����7�!�u�0�'�g������ƹ��E�����0�%�:�u��8����Cӕ��]��^�����w�_�u�!�%�?��������UF��X�����;��%�e�w�4��������A��d�����<� �0�>�2�}�ϭ�����V
��g��E���<�;�9�<�w�)����s�����X�����4�!�u�x�!�2��������9��^ ךU����0�!�u�w�8����Y����G��t��[���u�%�:�0�$�<����U����_��\GךU���0�<�_�u�w�}�ǿ�������Yd��U���u�&�0�!�%�����	��� ��D�U���u�0�&�3�%�.��������R��R-��\ʡ�0�_�u�u�w�}�%�������_��G��Hʦ�0�!�'��;�f�W���YӃ����=N��U���u�'�6�&�l�W�W��:����VF��RN�����&�3�'�!�2��6�������\��~�����;�:�;�u�9�}�'�����ƹ��T��]���&�!�u�4�'�8����Yӄ��ZǻN��ʴ�0�0�u�=�9�}�W���
����r��R��I���:�=�'�u�i�z�P��Y����_�������0�2�}�4�'�8��������9F�N��Xʖ�0�!�u�=�w�9����Y����G��C��ʶ�0�3�6�0�#�1����	ӄ��R��Y	��E���:�!�0�u�w�}�Z�������AF��C��ʦ�=�&��_�w�}�W�������P
��\(�����h�f�u�;�w�����������Yd��U���u�&�0�1�3�/����DӔ��Z��D>�����}�m�1�"�#�}�F��I���T������9�0��!�%�����P��ƹF�C�6���!�u�=�u�3�/�����Ƹ�VF��T��U���3�<�<�;�w�2�«�Y����W��PN�Eʡ�u�=�_�u�w�}�ZϷ�������DN��U���4�0�;�u�w�}�����Χ�E��[��3���:�u�u�u�9�}�%�������_�X�����'�9�6��4�2�W���Y����@4��C��6����%�|�!�2�W�W���Y�ƿ�V��S
�����h�'�&�/����������W	��C��D���e�u�u��$�����0����C ��C�����u�u�x�u�%�<�Ϫ�Ӈ��A����U���u�<�&�u�8�;�����Ơ�\��GN��U���;�u�=�u�9�8��ԜY���K��^������4�0�;�w�}�Wϻ�
���F�N�����1�'�&�u�j�/����Q����@��\����!�u�d�y�g�f�W���YӃ����=N��U���u�3�_�u�9�}����
��ƓF�'�����=�u�:�3�>�4��������$��zN��Cʾ�|�_�u�x��<�W���Y����U��R �����1�9�4�3�8�}��������9F��E�����4�%�0�9�~�}���������E�����1�0��8�;�������ƹF������!��!�i�w�����������^ �����&�0�1�1�%�.�^��Y�����V
�����!�<�0�i�w���������l�N��ʼ�n�u�0�1�'�2����s���F��R�����!�<�u�%�2�}�Fϼ�����V
�������u�:�3�<�>�3�W�������W��U������0�3�6�2�)�Jϭ�����@4��S*������%�}�`�3�*����L����F��X��1���4�i�u�<�9�9��������|��^��D���:�;�:�e�~�W�WϮ�����5��G�����u�7�2�;�w�}��������l��RF������>�u�=�9�}�W���T�Ɯ�C��Y�����'�6�<�;�;�-����ӕ��R��YN��U���!�<�u�<�2�}�ϩ��Ƹ�VF��E�����<�2�u�u�w�p�W�������\��C��U���&�;�0�&�#�}�Ͽ�
����WF��[�����'�0�u�:�>�;�Ϫ�Ӣ��^��T�����,�u�u�u�$�/��������c��N�U���;�1�r�r�q�.����0������Y��E���_�u�u�u��<����
����Z��R�����6��4�0�9�4���Y�����V�������%�g�k�}�1�������V/��^��N���u�u�&�'�4��������� F������=�&���'�o�}���Y���2��DN�����;�u�!�2�w�(�ϼ�Y���� �������7�!�0�;�#�8�5���Y����G��s=��M���9�6�_�u�w�}�4�������R6��R^��Hʦ�:�3��9�6�W�W���Y����Z��^ �����<�4�u�:�1�4����YӒ��^��_N��ʱ�9�4�1�9�.�}�W���
����U��R �����u�h�&�:�1�4����B���F��t�����0�!�<�0�w�`�W�������Z��g��E�ߊu�u�;�u�1�W�W���Y����V��=d��X���;�0�u�=�w�(���� Ӈ����N�����3�!�0�9�0�>����?����]F��^�����&�_�u�x�$�2����ӕ��X��^ ��U���u��a��4�0�������C��R��&���9��>�_�w�8��ԜY�ƥ���^ �����}�4�%�0�;�t����s���F�/��U���!�0�1�!�w�3��������V��C��ʼ�&�1�u�=�w��Cכ��Ƥ�_��^�����;�_�u�u�w���������]6��RZ��Hʦ�'�6��4�2�3����B���F��t�����!��%�d�k�}�4�������R6��R^�U���u�&�:�3�>�4����	���F��t�����0�!�<�0�l�}�W���T�Ə�V����U���!�%�,�u�w�}�������@%��Q�����<�0�u�u��<����
����Z��d��U���x�u�'�4�2�)�Ͽ����(��RN�����0�;�0�u�8�3��������\��X����� �7�'�_�w�}�W������A��M��8���y�g�u�u�$�2��������Z��H��E��e�e�e�e�g�m�G��I����F�=�[�ߊu�u�;�u�1�W�W���Y����V��=d��X���<�0�<�0�#�8�����ƣ�VF��E�����u��<�u�>�8����
������_��U���'�1�6�u�8�)��ԜY����V
�������u�=�&���e�W����ƭ�WF��RN��6ʑ��m�u�9�4�W�W�������R4��R�&���9��>�_�w�8��ԜY�ƥ���D�����_�u�u�u��8����5���F��C����u�e�|�_�w�}����Y����]��S	��&���9��>�u�?�3�W���Yӕ��V ��B����u�<�;�1�$�9�_������\F��G�U���0�1�<�n�w�8�Ϯ�����l�D-�����!�i�u��2�;��������]��c"�