-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����A��~ �����:��:�>�!�9�Z�������	F��_ �����8�;�x�u�%�:����)����P��g6��*��`�_�x��#�g�F������W��CחX���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�]�p�_���K����p	��E��ʛ�!�:�4�u�9�)�����Ə�A��V�����u�9�u�<�?�.�%�������K��V������&�'�8�9�.�>�������z��E�����x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��s����F��D�U���&�3�9�u�%�<�����Ƽ�\��D��U���6�u�:�u�?�}��������9K�N��U���u�<�!�'�8�<���Y����[��DN�����0�u��8�%�>��������@l�N��U���u�u�'�6��)��������GF��X��[���_�x�u�u�w�}�Wϊ��ơ�W�������4�;�"�6�;�(����Ӄ��A��^�����'��9��w�.����s���F�N��U���0�u�;�&�?�.�W���Y����R4��S/������3�0��{�4�W���Ӓ��]F��[�����!�0�x�u�w�}�W���Y����V��B��ʦ�6� ��!�x�}�����ƺ�_��@��U���6�8� ��;�9�������K�N��U���u��4�0�$�2����Ӑ��Z��E�����8�8�;�u��<��������@��C�����0�4�;�x�w�}�W���Y�ƺ�_��Q��R���0�6�:�>�6�)���� ����l�=C�U���u�u�u�&�6�<����0�ƥ�W��C�����=�'�u�&�9�*����Y����VF��D��U���:�!�0�8�:�/��ԑT���F�N��Uʓ�'�>�4�%�2��������J��s��'����1�0�&�1�.��������Z��V �����0�_�x�u�w�}�W�������GF��R
��ʼ�;�'�u�=�w�4��������@F����U���3�u�0�<�#�/�Lϊ��ƥ�9K�N��U���u�;�0�0�w�8����Y����w�������;�2�:�%�w�;����	����V��T��U���6�u�0�;�]�p�W���Y�����E�����6�;�7�u�"�5�Ϫ�Y����^��E��Yʰ�0�u�=�;�>�}�ϰ�ӟ����S�����x�u�u�u�w�}�W���Y����V��T�� ���<�;�u�4�>�}�3���+����W��D������u�4� �$�<����I���W�C��U���u�u�u�;�w�l�U�ԑT���F�N��U��x�u�&�u�?�}����ӂ��RH�r�����d�:�u�=�w�<�Ϩ�����R��=C�U���u�u�u�u�w�}�WϷ�����]��R�����"�0�u��#��!���Ӈ��V��@חX���u�u�u�u�w�m�W���,����[��R��ʻ�"�&�u�4�6�}�2������	��C�����u�4�<�u�6�<�}��Y���F�N��U���u�;�9�1�9�}��������[��D*�����4�<�u�&�2�)�^�ԑT���F�N��U��x�u�&�u�?�}����Y����@��V�����u�u�u�u�w�}�F���GӲ��@F�� ��U���4�<�u�3�$�)�}��Y���F�:��ʦ�2�4�u�&�#�0�W�������G	��s��#���1�;�_�x�z�}�W���Y���z��V��U���,�9�&�}��8��������w��NG��ʶ�9� �4�0�#�8��������]��C��U���u�u�u�3�2�}�$�������z��D������<�u�0�9�}��������C	��^ �����u�:�u�=�]�p�W���Y�����T�����u�0�1�u�8�/��������r%��Y��Mʶ�:�>�u�,�;�.�������F�N��Uʦ�!�'��9��}��������GF��\��Gʶ�6�0�u�:�1�:�����Ƹ�VF��P�����_�x�u�u�w�}�Wϳ�����A�������u�9�&�d�4�>�Ϫ�Y�������� ���1�!�u�'�:�0����U���F�N��Uʓ�'�!�<�u�2�.�ϭ�����e��SN��ʦ�4�4�0�1�3�/��������]F��RN�����1�x�u�u�w�}�W���Yۍ��G��[�����|�6�6�0�w�3����Y����_�CחX���u�u�u�u��}����Y����P��R��ʢ�<�0�4�1�#�8�W���ӂ��RF��X������u�4�4��0����U���F�N��Uʁ�u�4�6�u�?�}�4�������c��s��ʢ�u� �!�=�!�}����Y������D*�����<�0�z�_�z�}�W���Y�����T�����0�u�3�0�w�����������R��U���u�;�u�9�4�}����Y����Al�N��U���u�u��!��1����Y����c��b ��ʢ�9�u�0�4�w�5�W�������Z����U���9�u�:�6�2�)�}��Y���F���U���:�,�"�<�2�.����Uӕ��G�������<�0�4�<�9�9� ���Y����R/��^��Z���x�_�x�u�w�}�W���-����Z��^ �����,�!�'� �?�)����������^�����&�_�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T��Ɠ_��V�����y�"�'�n�w�(�Ϸ��ȿ�W9��P��D��{�9�n�u�"�8����W����A��D�����_�u�&�u�8�6�'�������Z��D*��[���n�u� �0� �/�Y���?����z��E����u� �0�"�%�s����	݇��l��Y��ʓ�4�!�;�0�'�/�����ƥ�9F��R �����u�u�>�4�'�8�'��� ����	F�������u�h�d�_�w�}�8�������u��X��U��<�u�;�0�2�}�J��s���X(��g�����;� �<�&�m�4�W�������	[�G�Uʥ�'�}�u�u�6�8����Y����\	��V �U����8�9��<�g��������T��=d��U���u�#�'�u�>�8��������PF��D�����u�0�u�<�#�/��������R�������;�&�=�&�y�}�Wϭ�����R
��N��U���9�4�n�u�w�.����Y����]F��V��¾�4�%�0��%�$���Y����G	�U��Xʀ�l�m�_�u�w�����/����\��YN�����;�_�u�u��)�%���8����@��Q��<���u�;� �&�0�8�E�������X5��G��%���,�9�x�u�8�3���B���fT�=N��U���!���%��g��������W��S�����|�u�x��o�l�W���
����z��G��Oʼ�u�<�;�1�f�}�������K�d_�D�ߊu�u��6�:�(�!�������F��X����u�u�&�6�"�����Y����w��x��¾�4�%�0��%�$���Y����G	�U��X���a�{�_�u�w��������	��*�����
�}��8�;�.���������Y��E���u�x�u�a�y�W��������]��G>�����6�n�_�'�?�)����Ӵ��	��q�����0�%�'�6�;�>�W���s�Ƹ�C��_��4���!�<�u�'�6�u�$�������A%��[��U���;�:�e�u�1�����ۍ��^6��T�����;�!�u�:�9�2�G��YӒ��VF��V�����<�u�'�4��<����Y����VF�N��U���<�;�1��%�$�ǵ�����P��^ �����u�:�;�:�g�f�WϪ�	�Ɵ�T��V�����<�u�'�4��3����Ӕ��T�	N�����<�;�1�a�w�2����I��ƹ��RN�����'�
�u�&�6�/�ǵ�����@6��t����1�"�!�u�~�2�W�������r��CF�� ���:�0�&�;��4�Ϻ�����O��N�����:�9�4��#�4�(���
Ӈ��R��d�����0��6�0�f�9� ���Y����UF��X�����!�'�>� ��2��������G��X����n�u�x�u�;�}��������Z��@�����u�=�u�4�2�9��������V�vN�����u�=�<�u�1�9����
Ӕ��F��Sd��X���:�%�:�4�6�8��������7��XN��ʻ�-�u��!������(�Ɵ�]��V�����u�<�;�9�6�.������ƹK�V�����u�;�<�0�6�:�����ƿ�R��R ��U���6�0�!�u�w�(��������G	��^�����!�0�%�'�]�}�ZϿ�
����V��N�����9�8�;�u�w�3��������7��DN�����:�1�<�0�#�8����Y����]Hǻ��ʜ��!��,�#�4�W�������`��[�����6�0�x�d�3�*����Y�ƣ�5��Y��M���4�
�}��:�/��������Z��S�����|�_�u�x�w�/��������^��V�����4�&�!�u�>�8��������\��X�����9�u�;�u�6�>�W���Y����JF��F�����!�u�;�!�2��������F��P ��U���!���9�3�4���;����R��T��]���!��9�1�2�<�W���Y����G	�UךU���;�9�&�'�8�4���=����A�������9�1�0�4�w�l��������\������h�u�:�=�%�}�I�������[�^��\��_�u�<�;�;�.����:����A�,������!�<�
�l�}�����ƿ�[��v��Oʅ�4�0�'�
�l�}�����ƿ�R��S/�����!�'�u�u�%�2����Q����C
��g�����x�u�:�;�8�m�L���
����_F��V������,�o��8�8��������l�D������!��,�w�}��������G]ǻ�����&�4�4�'��g�>�������l��N�����u��6�8�6�4�6���CӤ��_��z�����n�u�&�2�6�}�6�������\��T��4���!�_�u�<�9�1��������bF��v�����
�n�u�&�0�<�W�������G'��~N�4���8�'�
�n�w�.����Y����F��C/��$���6�8�'��f�}���T����X9��P���ߊu�x�=�:��4����s����]lǻC�6���!�u�u�0�6�8�W���
����\ ��s��<���9�1�!�u�6�>�W���Y����_���� ���8�;�u�;�#�8�'���,����l�G�����4�0�0�y��0�������Q��Yd��Uʼ�}��&�!�w�5����Y����w��~ �����<�0�i�u�8�5����GӀ��@�=N��U���<�u�<�<�0�8��������p
�������u�u�&�4�6�3����)����[��s��<���9�1�<�0�$�<��������Z��_��U��1�"�!�u�~�{��������_��=N��U���u�3�_�u�9�}����
��ƓF�C�����<�&�u�'�4�.��������G��DN�����;�4�<�u�2�<���� Ӎ��G��[�����u�,�9�&�]�}�W��7������C��#���1�<�0�4�3�.��������zI��V�����!�8�u�9�0�8�Y���Yӕ��G��[�����|�e�u�h�$�<��������Z��D*�����4�<��%�p�4���Y���F��V�����0�<�u�0�6�8�W���Oө��A%�������:�u�=�u��9�����Ƙ�Z��V�����=�u�'�6�9�)�W���T�ƾ�B��R�����0�6�;�?�$�}�����Ƹ��������'�6�&�<�0�(���Y����w��v��]���e�u�h�&�6�<������ƹF��s��4���}�|�e�u�j�.��������b]ǑN�����!��:� �>�� ��YӀ��5��~ ��ʼ�u��8�9�$�8�4�������\��XN����'�!�_�u�w�p�>�������VF��RN�����0�0�0�!�>�}��������G	��R�����3�'�!�%�8�8����Y����	��N��X���4�=��6�%�*� ���Y����G	��[��ʦ�2�4�&�4�3�>��������F
��X�����0�{�u�u�$�5���� ۵��z��OG��\��u��4�0��>����P���F��C��6����,��6�9�8�^��Y����`��C-���ߊu�u��6�:�/�>Ǎ�����KO�N�Uº�=�'�u�k�p�z�L���Yӕ��P��E��&���;�0�|�e�w�`�_������F�G����u�x��9�.�.��������W��D!�����;�!�u�0�#�)�ώ�����GF��G�����0�4�u�0�"�/����
���F��X���8�9��>�]�}�W������F�^�����2�0�2�}�6�-����PӒ��]l�N��Uʦ�'�:�<�0��>����P�Ƨ�R��V��1���,�x�d�1� �)�W���E�ƿ�A��^��&���;�0�|�u��)�!�������JF�N�����u�|�s�&�6�<��������@)��D���6�;�0�|�]�}�W����ƥ�l�N��ʥ�:�0�&�_�w�}�Zω��Ƨ�R��R�����9�u�&�d�#�8�3���Y����'��E��U���&�!�<�u�;�<���s���@"��V<�����&�!�'�}�'�����Q���F��E������6�;�0�~�6��������V
��C��\ʢ�0�u��8�;�.�������T��[��]���0�&�h�u�g�t�}���Yӡ��V��R>�����!�o�u�u�1�/�Ϸ�Y�Ƹ���Z>�����<�2�;�!�w�8�������F������u�'�6��#�/�'���,����F�N����>�2�>�4��.����Yۏ�l�N��Xǣ�:�>�4�&�#�/�4���0�ƿ�G��t��4����6�;�0�~�4�F�ԜY���K��X��ʦ�=�&��u��<����Q����]��F��D�ߊu�u�u�x�?�2�(���=����V��S
�����3�0��u��)�%���6����G'��=��<���-�}�x�|�w�}�W������l��d�����6� �u��6�)�����Ο�P/��R���ߊu�u�u�x�?�2�(���)����|��D>�����,��6�;�2�t��ԜY���K��X��ʦ�4�4�0�1�3�/��������F��s��'����3�0��.���������l�N��Xǣ�:�>�4�&�6�<�����ƿ�R��V��4���e�}�x�|�w�}�W������l��s��<���%��&�4�6�/�>��Q����9F�N��X���:�
�u��#��'���(ӕ��G��N?��\¼�d�_�u�u�w�p����&�ƿ�R��B�����&�4�4�4�>��Ǎ�����KO��d��U���x�#�:�>�6�.��������w��v��]����1�-�}�~�}�W���Tސ��\�������!�u��!��$�_���0����N��=N��U���x�=�:�
�w������ƿ�P��v��]����1�-�}�z�t�W���Y����[	��h��4���8�;�u��4�0����*����W����\���u�u�x�#�8�6�ϭ�����F��[����� ��9�1�%�u�������ZOǻN��U���=�:�
�u��>����5����@'��B�����%��1�-��t�W���Y����[	��h��4���8� ��9�w���������C��S��]���u�u�u�x�!�2����
����^)��~N������!�'���>����Pۏ�F�N����>�4�&�6�"�����8����|��E��&���;�0�|�<�]�}�W�������]��G>�����!�o�0�!�#�}����?����z��E�����<�u���]�}�W���Y����A��Z��]���u�u�u�u�<�<����)����P
��
P��&���9�&�0��4�8�W��Y���Z��P��O���_�u�u�u�w�}�8�������u��X��Kʾ�#�'�9�6��>���Y����]F��Y�����h�f�u�u�w�}�Wϵ�����G��RN��U��u�<�d�|�w�}�W���Y���F��N�����'�o�u�_�w�}�W�������R�=N��U���u�u��&�#�}�W���Y���F�N��H����&�!�u�w�}�W���Y���F�N��U���u�x�u�;�w�2����s���F�N������>�u�u�w�}�W���Y���F��Z��6���u�u�u�u�w�}�W���Y���F�C����&�1�9�2�w�}�W���Yӕ��R��V�����u�u�u�u�w�}�Iϭ�����R
��E�����1�-�}�x�~�}�W���Y����]F��X���ߊu�u�u�u�w��������F�N��U���u�h�u��6�8����	����V�^C�Y���u�u�u�u�z�}��������Vl�N��U���&�!�'��;�����Y���F�S����'��9��.���������J�N��U���x�:�!�7�8�8����Y���F��g�����u�u�u�u�w�}�W���Y����c��R/��]����1�-�}�~�}�W���Y���F���U���<�;�_�u�w�}�W���=����]0��^
��U���u�u�u�u�j�}�3���/����r��G��X���u�u�u�u�w�}�W��Y���Q	��R��U���u�u�u�&�6�<��������@)��D�����k�&�4�4�3�9��������`��Y
��\¼�d�y�u�x�>�}������ƹF�N��U���!���%��}�W���Y���F������,�}�|�<�f�q�W���Y���F�N��X���;�u�<�;�3�W�W���Y���@"��V'�����u�u�u�u�w�}�W��Y����R'��fF�]���|�u�u�u�w�}�W���Y���F��N�����}�u�u�u�w�}��������R
��N��U���u�u�u�k�$�<��������5��~ �����|�u�u�u�w�}�Zϱ�ӄ��_��=N��U���u�u��!��<�6�������U��x��H����!����;���� ۵��z��OG��\���u�x�u� �w�3����s���F�N����� ��u�u�w�}�W���Y���F��V������6�;�0�~�4�[���Y���F�C����&�2�0�}�w�}�W���Yӕ��G��C?��U���u�u�u�u�w�}�Iϭ�����J7��G�����}�|�u�u�w�}�W���Y����F��^	���ߊu�u�u�u�w��������F�N��U���u�h�u��4�0����*����W����\���u�u�u�u�z�}��������l�N��U���&�6� ���}�W���Y���F�S���� ��,�}�'�����Q����F�N��U���x�<�u�&�0�8�_���Y���F��v������9�u�u�w�}�W���Y����r��Z/��<�6�;�0�|�>�q�W���Y���F���U���;�1�_�u�w�}�W���8����|��T��U���u�u�u�u�j�}�6�������5��~ �����|�u�u�u�w�}�W��Y����@��R
��U���u�u�u�&�4�(�8�������F�N��U���k�&�6� ��1����Q����]��F��Y���u�u�u�x�8�)������ƹF�N��U���6�8� ��w�}�W���Y���F������ ��,�}�'�����Q���F�N��X��� �u�<�;�3�W�W���Y���@'��B�����u�u�u�u�w�}�W��Y����F��C/��$�6�;�0�|�>�t�W���Y���F��CN�����}�u�u�0�3�:�����Ƌ�]��C�����<�&�_�u�w�.����6����`��Y
��\��u��6�8�"�����	����V�\ ��%���0�&�;� �>�.�_������\F��d��Uʦ�6� ��!��-�>��������T�� ���,�}�%��3�%�_�������V��Y	�����}�`�1�"�#�}�^�ԶY�Ʃ�WF��Y�����0�0�4�0�%�>��������9F�C�����=�u�'�6�$�4�ϫ��ƾ�D��V�����&�8�u�4�6�-��������9F�C��ʻ�0�u�;�,�8�8��������e��SB��ʶ�;� �0�4�.�}�ϩ��ƹ�VF��RN�����:�0�_�u�$�>��������WF������4�<��,�g�u�9�������@��b ����_�;�u��l�