-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����A��~ �����:� �<�{�?�W�Zϟ�����,��YN�����4�u�;�u�8�8�4�����ƴF��^	�����'�?�6�o���(��L���"��RT��Bʟ�9�u�e�d�z�W�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K��C�����e�d��%�%�:�ϐ�����_F��D�����&��'�:�6�4���Y����a��C�����#�1�x�u�6�4����0����F��C�����;�9��3�%�<����T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C����x�u� �%�$�g�W���
Ӌ��F
��T�����:�0�%�:�2�.��������\��_�����<�;�9�x�w�}�W���Y�ƥ�G��X�����x�_�x�u�w�}�W���-����^	��[�����&�4�;�"�4�1��������E����ʦ�!�'��9��W�Z���Y���F��D�����u�!�"�9�w�<�����Ƨ�E��[��3���:�u�:�3�>�4��������9K�N��U���u�:�3�:�w�����Ӈ����C��ʡ�0�u�<�=�#�8��������W��
��ʼ�u�=�_�x�w�}�W���Yӕ��U��R	�����{�x�_�x�w�}�W���YӲ����T����� �<�u�<�;�<�Ͽ�Ӊ��G��Z�����u� �%�!�w�2�Z���Y���F�D/�� �����!�u�%�<�Ϫ�ӕ��P��B��$ʺ�!� �u�=�#�4�W������F�N��U���=�;�&�6�"������ƭ�@��D@��;���1�!�u�&�$�4��������G��D�����u�u�u�u�w�}��������Q��D�����u��!���1�ϩ��ƺ�_��S��U���u�,�9�&�z�}�W���Y���_��EN��U���!���%���}��T���F�N�����4�4�<��w�3�����ƥ���E��ʻ�"�1�!�u�8�?�W�������]��C�����'�0�_�x�z�}�W���Y���u	��\=������'�,�9�w�}�[ϭ�����R��S�����&�!�;�6�9�<����ӏ��V��=C�U���u�u�u�:�1�8�W���Ӓ��Z��E�����<�&�u�4�'�8�W�������[�������'�n��<�w�.�Z���Y���F�Y�����0�4�&�u�2�}����������P�����3�>�4�%�2���������[�����߇x�u�u�u�w�}����ӂ��RF��YN��U���=�1�!�u�?�}�������V����ʼ�u�&�;�!�.�)�����ƪ�Al�N��U���u�u�=�u�"�/��������R��Y@�����u��!��6�����
����V���� ���4�0�w�e�{��F�ԑT���F�N�����d�w�_�x�w�}�W���Y���F�;��U���u�0�0�!�3�)�Y�������GF��X�����4�!�#�9�3�9���T���F�N��U���u�u�<�6�"�4�ϰ�ӂ��RF��R ��1�����9�1�6�.����W���F�N��U���e�u�k� �2�)�ϭ�����]��D�����u��0�0�#�m�����Ơ�@��V��U���4�_�x�u�w�}�W���Y���F��Y�����u�0�u�4�6�*����=����]0��^
�����!�|�_�x�w�}�W���Y���F�;��U���u�=�'�u�2�8�Ϻ���ƴF�N��U���u�d�u�k��4�W���������^
�����!�_�x�x�w�}�W���Y�ƛ�V��R�����<�u� �=�3�)�W���Y������C�����u�<�0�4�9�*��������\ǶN��U���u�u�&�4�#�}��������GF��C�����=�u�4�!�3�)�W���ӑ��_F�������u�:�!�0���}��Y���F������3�9�:�<�0�6��������p��RN�����{�x�_�x�w�}�W���YӲ��@F��P ��U���!�8�u�9�0�8�W���
����e��S'�����x�u�u�u�w�}�W���Y����GF��P ��ʴ�0�0�%�6�2�}�϶��ƨ�U ��R �����9�;�u�0�6�.�}��Y���F�:��U���9�"�;�u�6�<����
ӂ��P��RN��ʧ�$�<�0�0�#�;�ϻ��ƿ�T��d����u�u�u�u�w��W�������P��R�����3��9��'�����Y����R
��[��U���u�:�3�<�>�3���Y���F�N�����&�!�'��;��W�������2��DN�����!�0�6�'�2�-����ӂ��RF��EN�����u�u�u�u�w�}��������]F��R
�����0�6�u�=�w��W�������_	��DN�����u�3�0�_�z�}�W���Y����`��C-�����4�&�'�&�w�)����
����J��DN��U��� �0�:�!�#�8����ӂ��Rl�N��U���u�u�0�:�.�/��������@F��B��U���9�u�:�'�6�}����������VN�����0�:�,�_�z�p�W���Y���F��V�����<�u�;�u��)�%���8����@��Q��<���=� �1�x�w�}�W���Y�ƫ�GF����ʠ�<�u�u�>�6�<����=����F��T��U���0�u��4�#�<����s��ƴF�N��U����u�4�0�w�*�W�������\F��^�����!�0�u�0�3�9��������[��e"������8�'�0�{�p�W���Y���F�������=�u��0�1�<��������JF��V�����0�z�u� �#�5��������W��=C�U���u�u�u�c�4�2���� ������R��&���!�4�6�;�6�.��������]��[��U���9�u�3�0�]�p�W���Y�����C�����;�_�x�x�w�}�W���Y�ƿ�G��t��:���u��4�0�"�q��������R
��N�����0�1�1�'�$�����6����]ǶN��U���u�u�&�4�6�(�'���0ܷ��A��[�����<�0�u�0�$�2�ϱ�Y����P	��R�����2�<�%�!�z�}�W���Y���@��V�����u�=� �1�5�}�����Ƹ�VF��O�����&�<�2� �>�s�W���
�ƿ�T��Dd�U���u�u�u�u�%�}�����Ʈ�-��R�����4�!�'�6�4�8�W�������]��X�����6� � �4�>�3���� ���F�N��Uʺ�u�=�u��w�3��������r%��^�����0�&�=�&�w�2�W�������P��T��U���9�&�4�1�z�}�W���Y���R��Z�����9�u�=�u�%�9����W���K�N��U���u��6�;�#�3�Ϻ�����]��@��ʶ�0�3�6�0�#�}����
����JF��^חX���u�u�u�u�>�.����W�ƚ�_��A�����4�2�u�'�:�m����7����\��D�� ���&�x�d�_�z�}�W���Y����~��Y�����<�u�9�:�"�8�W�������_����U���'�6�u�0�3�<����
Ӏ��9K�N��U���u�!�0���.�W���Ӓ����E��U���4�<�u� �#�-��������Z��T�����;�<�2�x�w�}�W���Y�Ư�V ��T�����_�x�u�u�w�}�Wϊ�Ӏ��_F��G�����0�4�u�=�8�:�W���
Ӌ��F
��^��%��� �<��6�:�8��ԑT���F�N�����&�_�x�u�w�}�W�������f��c�����4�u�h�>�8�;�4���)����V
��E��8���<�0�0�4�w�}�'���,����P��s���߇x�u�u�u�w�}�W���Y���F�N��U���h�d�u�u��8��������\�CחX���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�]�1���� ӏ��VJ��X�����&�u�0�0�$�9��������H��[UךU���u�0�0�;�:�/����݇��l�B�����{�>�� �>�4����
�ȭ�_]ǻ��U���>��2�&�y�1�L�������\��g������!�'�{�;�f�}��
����V�������!�
�3�_�>�/��������p	��{�����'�'�u����}���Y����z+��T�����!�{��n�z�}��������G��D�����_�0�!�!�w�/��������A	��Y���ߊu�0�0�<��}�Wϵ�����@6��t����<�u�;�0�2�}�J��s���X)��E�����6�:�u�u�9�4������� ]ǻN��8���;�!�;�0�m�4�������O��N�����u�u�4�0�2�}�W�������R��N��&���9��>�o�>�}��������9l�N������9��u�w�3��������F�D>�����u�o�<�u�9�4��������V*��P��X��1�"�!�u�~�}�Zϋ�@��ƓF�D=�����9��!�o�8�)��������F�D>�����!�o�:�!�"�.����Q����@��Y	��U���u�:�;�:�g�f�Z���K����9F�C�!���3�9�:�<�0�.����
ӕ��F
��U�����0�u�u�,�;�.� ���Y����V��N��X���:�&�!�'��1�>�ԜY�ƿ�R��Y8�����u�;�7�:�2�3�}���Y����R4��S/������3�0��w�}�ϫ�
����WN��S�����|�u�x� �y�W�W���Tӕ��G��g��<ń�&�:�9�u�8�)��������W����U���6�_�u�u�z�>����Y����AF��C��6����u�&�0�#�s�W���
����z��G��Oʼ�u�<�;�1�f�}�������K�d_�D���u�&�4�4�9�4����Y����Z��SF�U���;�:�e�n�z�}�F���s�����C�����<�u�u� �w�2����B�����C�����1�0�&�3�$�)����Y����F��P ��]���:�;�:�e�l�p�W��K�����C�����u� �u�<�9�9�F�������V�C�&��d�u�u�&�6�<����CӉ����Y��D���:�;�:�e�l�p�W��W��ƹF��v�����u�u�;�&�0�8�_������\F��N��Xʆ�c�b�u�u�$�>����(����]F��P ��]��1�"�!�u�~�}�Z���M����9F�C���� ��!�6�������ƣ�_��RN�����!�1�!�u��>����V���F������u�:�0�3�%�}�W���Mˣ��]��E�����1�1�!�u�8�)�W�ԜY�����P��ʑ��m�u�:�'�3���Y����r��Z!��9���u�u� �u�>�3���Y����G	�U��X���a�{�_�u�w���������bF��X�����0�}�b�1� �)�W���Y���`R��dךU����6�8� ��1�������\	��V �U���&�6� ��#�}�W���Y����V� N�����u�|�u�x�w�i�Y�ԜY�ƿ�P��x��U��� �u�<�;�3�i�W������O��C�&��l�0�1��6�)����	����f��d�����!�6� �0����������]��G>�����!�<�_�u�4�0����ӵ��pU��=N��U���!�}�u�u�w�>����ƿ�W9��P��O���e�n�u�u�w�9�MϷ�Y����_	��TN�U��n�u�u�u�4�}�W���
����\��T��R��_�u�u�u�w�}�ϭ�����Z��R����1�"�!�u�~�W�W���Y����\��D�����6�_�u�u�w�n�W����ƿ�W9��P��N���0�1�6�8�8�8��ԶYӕ��]��D=��'����1�0�&�w�}���������Y��E�ߊu�u�u�u�w�}�W���Y���F�S�����'�u�k�r�p�f�Wϭ�����@5��e��4���0�&��u�m�.��������V��EF����!�u�|�_�w�p�#���*����W��D��@ʷ�!�|�=�&�6�0����Ӑ��F��QN�[ʂ�u�4�0�!�w�<�ϭ����K��RN��ʻ�#�'�2�<�0�)�W���Y����P��DN�����0�u�1�'�$�s�W��Y����^��Z��&���4�1�0�&�"�8�W�������^��SN��U���u�:�9�"�9�}��������F���]���9�0��!��1��������P
��\(�����~�8�-�&�6�<��������@)��D�����u�_�u�x��%��������r��R�����!�;�#�9�3�4�W��Y���~��A��ʾ�<�!�'�4�6�8����
����U	����6���b�3�'�f�w��}���Tӫ����[<�����'�&�u�:�w�%�8���
����F�N��G���d�h�f�_�w�p�:���
����V��S
�����:�u�-��w�.�W��Y����F��N�H��{�u�&�2�6�}�3���6����^��N�����2�6�#�6�8�u�@Ϻ�����O��N�����u��!��#�2����Y����_	��T1�����}�b�1�"�#�}�^�ԜY����R
��s��8��� ��o�&�0�8�_������\F��T��]���0�&�h�u�g�t�}���������C������o�&�2�2�u�@Ϻ�����O�
N�����&�h�u�e�~�W�W��Y����WF��R������6�:�&�1�/����Y����_��E��X����=�'�#�;�8�W���ӈ��9F�N�����0�!�1�u�1�$����������RN�����0�0�!�'�;�)�����Ƹ�Z��X
��U���u�0�1�u�?�3����ӕ��C	�������x��u� �'�/�W���6����_	��q�����3�d�!�0���Dݛ�����]���� ���;�!�7�_�w�p����Y����P��A��U���!��!�0�6�}����Y����_F��X��[���&�7�,�0����������]��CN��U���0�0�u�4�0�}�W������l�C�����,�>�#�'�;�>�1����ƥ���E��ʱ�3�;�1�7�w�+��������R��h�U���u�=�&�4�4�4�����ƣ�_��B�����&�6�u�4�0�s�WϽ�����GF��R�����9��6�:�w�}����?����A4��P�����u�u�u�u�w�}�W���Y���F�N�U���0�6�:�>�6�)��ԶY���e��SN��6ʳ�'�!�<�u�8�(�Ͽ����F��_�����0�u�4�0�9�)����s�����C�����4�0�;�!�$�-�������K��XN�����!�2�0�!�%�+����Y����w��=��U��� �!�'�u�2�9�W�������VHǻ�����u�%��;�2�)��������AF��Y	��Gʱ�"�!�u�n�w�p�W�������|��T�����!�'�<�u�9�/��������V��NN�����2�
�{�u�z�}��������G��B�����u� �%�'�$�.��������9F��X �����>�0�<�,�'�����Cӵ��a��R1��O����8�9�&�2�����s����\��V ������%��9�.�}�W���Cӏ��V��T��F�ߊu�:�&�4�#�6��������P��R��U���;�0�0�u�j�6��������R��EN�D�ߊu�:�&�4�#�6��������G��R��U���;�0�0�u�j�}��������P6��R*���ߊu�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�v����)����V
��=N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�~�>�%�>��������V
��dךU���;�9�&�!�%��������	F��X�����!�'�>�'�4�3��������R�_�����:�e�_�u�w�}�W���Y���F�N��U��u�:�=�'�w�c������ƹ��Y�����&��9�,�w�}�W�������GN��A������6�:�u�w�}�������F�N��U���u�u�u�u�w�}�W��Yۉ��V��
P�����'�u�k�r�p�t�}���������C�����0�4�u�o��2����������R�����4�!�'�x�f�9� ���Y��ƹF�N��U���u�u�u�u�w�}�W��Q����A�	N�����n�u�&�2�6�}�3���+����U ��C*�����o� �&�2�2�o����&�Χ�E��[��3���:�u�u�u�8�3���s���F�N��U���u�u�u�u�w�g�WǱ�����X�X�����k�r�r�|�]�}����ӕ��G��R��U���2�0�d��/��������P
��\(�����x�d�1�"�#�}�^���Y���F�N��U���u�u�u�u�j�u����
���	��R��H���e�|�n�u�$�:����=����w��NN��U���;�1�m�'�6��_�������P��T��U���u�:�;�:�g�W�W���Y���F�N��U���u�u�o�u�8�5����G�Σ�[��S�R��|�_�u�x�w�<�ώ�����Z��Y�����<�&�1�3�2�8�Ͻ�����Z��DB�����4�=�6�0�1�>����Y���R�������,�1�1�!�{�.����
Ӓ����B�����;���3�;�8�YϜ�Y����TF��N�U���3�'�;�u��1��������R��YN�����'�6�&�<�0�3�ϩ�Y����[F��T�����<�<�;�_�w�p� ���Y����A��CN�����<�u�=�u�6�<�}�������]��q�����!��9�,�m�4�������X)��E-�����6�:�u�u��>��������9F�N�����4��1�0�$�4�W�������V��E�����#�9�0�{��}����Ӊ������ʷ�!�_�u�x� �}��������[��X �����4�!�%�'�w�8����
����R��C�����!�;�u�4�#�;�������K��V�� ���'��1�0�$�W�W��?����G��Z��&���4�1�0�&�6�<����Y����R��[����� �4�0�!�2�0�������F��V�����1�'�&��1�8�Y���T�ơ�KN��V�����1�'�&��1�8�^������w��e��4���0�&�3�&�#�3�W���?����A"��V*���ߊu�x�:�_�w�p����
����a��v
�����3�&�!�u�w���������P��E������!��4��9��������z�N�U���u��!��6�����
����V������:�>�4�!�%�v�F���
����_F��V�����1�'�&��1�8�W�������V��X	�����}��0��8�6�������F��@ ��U���u�u�u�u�w�}�W���Y���F�N��U���h�}�!�0�$�`�W��P��ƹ��Y�����3��!�u�>�3���Y����G	�UװU���u�<�<�u�?�}�����ˣ�GF����U���;�9�u�=�#�<�Ϲ�����\F����ʼ�u�4�,�u�z�}����
ӄ��R����ʴ�3�6�u�;�>�8����Y����@Hǻ�����!�u�4�
�6�2��������l�V�����0�8�-�3�9�(�W���
����V��S
�����u�<�;�9�>�}�N��YӇ��A��C�����4�:�!�:�w���������_��N�����u�&�w�w�]�}�Z¨�����Z��V��U���#�:�>�&�0�3�}����ƓF�-�����!�0��4�2�<�Ϛ��ƨ�_��E�����&�u�x�u�?�}�����ƣ���DN�����0�&�;�u�8�)�ϰ��Ƽ�\��D��U���!�_�u�'�4�.�_���	����XOǻ���ߊu�u�3�'�$�3�(���۵��C
��[�����_�u�u�u��<�������Z������0�4�}��6�8����^����W��X����u�u��4�2�3�}���Y�ƿ�R��R�����!�0�4�u�j�}�3���+����U ��C*������!��4��;��������Z��N�����u�|�s�&�6�<��������@)��D���ߊu�u�u��#�����Y���@"��V'�����&�4�4��;�$����T�ƨ�D��^��Sʦ�4�4�;�<�2�f�W���Yӕ��G��R��U��u��!��2�<�_�������_��_��X���:�;�:�e�w�}�3���0����V7��N�����<�n�u�0�3�-����
��ƹ��C�����1�0�&�3�$�)����D�ƿ�R��R�����!�0�4�}��8��������\�_�����!��!�w�`��������R��x�����>�4�!�'�z�l�L���
����|��R�����4��9�,�<�+��������G	��N�N���&�=�&��#�a�W�������_��\!�����6��6�:�w�}�^�ԶY���g��Z�����#�9�1�&�6�<��������@)��D��ʼ�u�{��:�#�.����������C��U���;�!�!� �y�}�Z��� ����@��C�����0�:�3�u�6�.����=����V��S
�����3�0��u�j�o�W�������GF��s��'����1�0�&�1�.�����ƥ�E��SB��ʸ�,�2�;�'�#�}�Ϸ�����5�������u�2�0�!�%�)����H���@��E��U���:�n�u�x�w�$�����Ƹ�R��V���ߠu�x�u�'�6�8����*����%��T�����u�0�4�u�2�4����s���'��^ �����<�!�u�4�"�}�Ϫ��ƨ�_��^�����!�u�=�u��}�Ϭ�
������DN�����9�!�'�u�'�2��������GJ��Z��6���_�u�0�<�]�}�W�������GO��_��U���u�&�!�'��1�3��� ���	��R��H���4�&�|�_�w�}����Y����]��S	��&���9��>�u�?�3�W���Yӕ��R��V�����u�h�u��6�)��������@5��E�����9�,�=�2�z�}�������F��C��6����n�u�u�2�9���YӃ����T��N���x�u�;�<�#�/�����ƺ�_��X�����1�9�,�6�6�3����
����\F��V�����;�-�u�'�4�.������ƹK�T�� ���<�;�u�=�$�9��������V��_�����4�1��4�2�9����W����`��C-�����u�h�u��6�)��������X)��E�����6�:�u�u�~�W�W��Y����G��_������9�1�1�;�$����
����9F��E������&�!��:�1�4���s�Ʈ�T��N������&�!�u�?�3�W���Yӕ��G��[�����u�h�}�!�2�.�J�������l�N�����'�&�;�
�3�8�$�������F��R ךU���u��!��;�9����Y����w��a�����4�}��!��1��������T�
�����e�u�u��#��!������F��SN��N���0�1�%�:�2�.�}���Tӧ��Z��E�����u�4� �u�1�)��������P��YN�����0�&�;�u�8�)�ϰ��Ƽ�\��D��U���!�_�u��#����������C�����0�4�}��2�>��������K�UװU���u�'�4�0�#�8��������r��R�����!�� �!�%�}�Z�������@F��R
��ʦ�9�6�u�=�4�}��������G��S��U���3�u�0�<�#�/�W���Y������C��8���{�_�u�x�v��9���Y����g3�������4��1�0�$�;��������GF��V ��U���0�<�!�9�w�;����+����9F�N�����'�&�7�6�"�8��������P/��E�����:�3�9�0�6�9����
Ӏ��@��X�����4�_�u�x�4�2�Ͻ�����R ��EN�����u�0�&�0�#�2�Y���	����@��V�����|�u�7�2�9�W�W���Ӕ��Z��R
��]���%�0�9�|�#�8�}���Y����VF��RN��9���:�&�:�0�#�8�3���Wӵ��@F��RN�����u�:�u�"�w�8����WӠ��@��RN��ʧ� �0�u�u�z�}��������R��R��ʡ�8�u��4�#�<��������G��NN�����;�u�:�!�2�/��������@�N��X���0�:�1�u�9�)�Ͻ�����D��RN������9��u�$�1� ϩ�Y������E��U���u�0�!�&�:�1����Y���Z��R�����u�:�1�u�?�.� ����ƿ�^�������!�:�0�3�8�}��������W��D�����u�x�u� �?�<����
����VF��SN�����=�u�4�0�6�9����s���K��_��4���-�0�!�u��8��������\��V�����!�0�:�1�$�}�Ϫ��ƣ���������4�!�4�4�3�W���T�ƭ�@��DB��ʾ�#�'�9�6��>���Y����V��^�����9�&�4�!�%�)�ϸ�����]�N��X���=�'�3�'�w�;��������R��Y�����&�4�'�4�.�.����Y����[��e"����3�'�!�0�2�8����Y���G��z/�����u�&�u�&�$�2����Ӈ��A�������4��1�0�$�;��������|��t�����!�'�x�d�w�}�Z���Ӓ��	��R�����u�3�;�"�$�0��������V�������!�u�=�u��}�Ϫ�ӕ��VF��Z�U���x�u��!��<�6�������U��~ �����u�;�4�?�$�0����Ӈ��\����U���u�4�%�0�w�5�Ͽ����K�Y�����=�u�0�:�.�$�����Ƣ�^�������9�&�w�0�3�3�UϷ�Y����C
��g�����u�u�{�u�w�p�W���Y����GF��R��ʡ�0���"�;�}����
ӕ��A��^ ךU���x�&�4�4�2�9����
����@��YN�����'�9�6��4�2�W���Y����`��[�����6�0�x�d�y�}�W��Y����w��e��4���0�&�3�&�#�3�\ϵ�����\��V�����>�4�%�0��/����s���K�`��U���0�u�4�6�;�)����������Y��U���'�4�u�=�w�4��������GF��RN��6ʢ�9�u�&�{�w�}�Z�������[��^��U���8�;�u�&�#�8����
�ƨ�G��V���ߊu�u�u�3�$�)��������R��t�����6�<�0�0�6�p�^Ϫ����F�N�U���;�"�u�'�w�2�W�������]��S��U���u�0�0�!�$�0����
ӕ��A��^ �����&�u�{�u�w�}�W��Y����_�������u�=�u��w�4�ϫ�ӏ��@��R
��ʦ�4�4�0�1�3�/��������]l�N��U���u�=�'�3�%�}��������V
��R �������0�%�4�.����������V
�����u�u�u�u�z�}�3���+����W��D������u�u��2�>��������K�d��U���u�<�u�:�w�����/������Yd��U���u�u�&�4�6�8��������U ��CN�U���!��4��3�8����
����M��x�����>�4�!�'�z�l�}���Y���K�`��U���&�4�!�"�>�4�Ϻ��ƥ�G	��_��'���;�u�,�9�w�8�����ƿ�R��E�����u�=�u�0�2�)�W���Y���F��Z��U���9�7�u�'�#�8�W�������a*����U���9�&�4�!�%�*�W���Ӓ�� ��D�����;�_�u�u�w�}�Zϸ�Ӓ��+��d��U���u�x�u��#��!���Ӂ��@F����ʰ�!�!�u�;�w�$����������C��%�����u�:� �}��ԜY���F���ʳ�'�!�0���*����Y������E��U���u�<�&�u�;�0�����Ƹ�VF��tN��&���9�&�0��4�8�Z��s���F�C�����0�u�'�u�8�}����Ӓ��5��N��ʇ�4�u�1�'�$�}����Y����G��=N��U���u�9�0�u�w�}�W���
����a��v
�����3�&�!�i�w���������A��x�����u�u��0�4�2���������Z������6�0�_�w�}�W����ƥ�lǻN��Xʜ�u�u�0�u�6�>�����ƥ��������2�!�<�u�.�1�[Ϫ�ӫ����R��U���u�0�!�1�#�W�W���TӃ��^���������u�3� �}��������R��^ ��U���u��u�=�$�>����Y����`��@�����u�x�!�>�w�<�ϱ�Y����]��R
�����<�2�u�3� �}�����Ƽ�@��PN��ʱ�!�y�"�u�?�;�W���s���K��S
�����:�'�4�u�?�}��������]��YN��ʆ��_�u�u�z�����Ӎ��CF��V�����1�'�&��1�8�W���Iӑ��]F��R�����:�0�!�8�w�4����Y����P��B�����_�u�u�x�5�4�ϵ�����\ �c��U��� �0� �u�?�3� �������@"��V<�����'�&��3�2�}�ϼ�Y����Z��N��X���'�0�,�u�>�8�W�����ƹF������:�u��!����������w��e��4���0�&�3�&�#�r�W�����ƹF�N��U���!��4��3�8����
���F��V�����1�'�&��1�8�W���B���F��Y
���ߠu�u�u�x�w�4��������a*��S
�����4�6�9�!�8�}�Ͽ�����G��Q�����0�4�u�;�w�2����Y���K�Q��U���u�:�`�7�#�s�W���Yӕ��_4��S/�����u�h�u��;�8�3���=����9F�N��U���u�u�u�u�w�}�W���������C�����1�0�&�3�$�)����+����W��D�����=�n�u�u�2�9���s�Ʃ�WF��X���ߠu�x�u�'�6�8��������^��E��'���0�1�4�1�2�.�Wϭ�����W'��E��&���i�u�!�
�8�4�(�������`��R�����&�|�_�u�z�}��������[��fN�����0�:�<�&�w�	��������^��Z�����<�=���w�2����Y����F��D@ךU�����o�u�1�/�>Ϸ�Y�Ƹ�W��P�����_�u�u�x�?�2�W���:�ԉ�5��t]��<���u�x�#�:�<�<����*����V%��=N��U���=�:�
�u�w�}�3���0����V/��d��U���#�:�>�4�4�}��������Z��s��#���1�0�4�}��)�>���=����K��s��#���1�0�4�u�w�t�}���Y�˺�\	��VN��Uʦ�'��4��3�8����s���K��X��ʤ�u�&�4�4�"�����0���F�A�����$�d�:�0�]�}�W���:�ԉ�	F��{-�0���u�u�%�'�w�<�W�ԜY���F��\N��U���%�0�9�y�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���x�u�;�u�w�}�WϺ�Y���@"��V'�����}�|�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N�����u�u�u�0�w�c��������Z��s��#���1�0�4�}��)�>���=����K��s��#���1�0�4�u�w�t�[���Tӏ��F�N�����h�u��9�2�9����
����F�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�x�w�3�W���Y����F�	N����� ��8���q�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���:�_�u�u�w�}�D���GӉ��]O��N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���K��BdךU���x�=�:�u���E���*����#��N��Xǣ�:�>�4�6�<�����:��ƹF������u�u�u��#��'���(ۯ�F�C�����4�6�u�!��)����ە��G��[�����}��!�������TӍ��G��[�����u�u�|�_�w�}�Z�������RF�D=��'����1�0�&��W�W���T����X9��FN�����4� ��8���}���Y�˺�\	��VN��Dʺ�0�_�u�u���E���Y���� T��N��Uʥ�'�u�4�u�]�}�W���Y����X��V�����y�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N�U���u�u�u�u�3�}�J���=����]6��R?��\���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���ZǻN��U���0�u�k�!��)����ە��G��[�����}��!�������TӍ��G��[�����u�u�|�y�w�p��ԜY���F��N��U���9�0�1�1�%�.�$���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���x�u�;�u�w�}�Wϯ�Y���@"��V!��6�����y�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N�����u�u�u�f�w�c����P���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���TӉ��F��SN�����!�u�0���f�}���TӶ��V
��RN��ʆ��:�!� �$�)�W�������G��Y	ךU���6�&�}�4�'�8����Yӄ��ZǻN��ʧ�&�;�
�1�2�����:���G��=N��U����!��8�"��K���������C�����7�|�_�u�w�}�3���4����G7�
N�����}��!��#�2����s���V��^�Uʰ�1�%�:�0�$�W�W��Y����G��_�����<�<�;�u�6�>�����Ʈ�\��N����>�0��4�#�3��������R
��N����>�4�&�0�#�/�4���Y����A��[�����x�=�:�
�w������ƿ�\��x��G���:�;�:�g�]�}����0����C%��Q�����u�;�<�,� �/�Y�������V��X��6���u���_�w�}�����ơ�CF�N��Uʾ�#�'�9�6��>����GӍ��V��X�����'�u�x�u�9�}��������UǻN��U���6�;�!�;�2�}�W��Y����z��V ��\���u�u�x�<�w�4���������CN�����u�u�u�4�2�8�W���Y�����D��U���u�u�u�u�w�}�W��Y���Q	��R��U���u��8�9��6�W���Gӵ��C
��[�U���u�u�u�u�w�p�W���Y����_	��Td��U���&�0�!�'��1�W���
����G%��T'��U���u�u�u�u�z�}��������]l�N�����&��u�u�w�c����
����F�N��U���u�u�x�u�9�}�������F��@ ��U���u�u�u�&�8�;�8���Y�����R�� ���g�1�"�!�w�t�L��Y����@��R
��Eʱ�"�!�u�|�]�}�4�������F��@ ��U���i�u�:�=�%�}�I���^��ƓF�-�����!�0����}�Z¨����� ��T�����9�'�4�u�6��W������l��q�����=�<�u��4�3������ƹK��_��*����&�4�!�6�>��������P"��V��6���3�4�6�<�2�8����Y��ƹK��_��*����!��9�3�)��ԜY�˺�\	��VN������u��0�1�(�}���T����X9��D*�����&�4�4�0��)�}���T����X9��D/�� ���u��6�8�9�W�W�������RF��T��:���6�u��6�:�(�;���s���E��\1����� ��!�&�4�(�8���s�Ɓ�P/��R �����:�>��4�#�8��������N��{GךU���0�0�<�u�6�}�}���Y�Ƨ�Z��~ �����h�u��6�9�)����I���F��N�����;�u�u�%�%�}����s���F��Z��6���u�u�k��:�1�4���Y���F�N��U���u�u�u�u�w�}�W���T�ƥ�F��S1�����u�u�u�&�6�<����Y�����RB��U���u�u�u�u�w�}�W���Y���F�N��U���x�<�u�7�8�8����Y����a��V�����h�u��4�#�<�����Χ�\��t��%����9�,�x�f�q�W������\	��V ךU���u��!��w�}�W��Y����R+��x��Y���u�u�u�u�w�}�W���Y���F�N�U���u�<�;�1�f�}�������F�D-�����u�u�u�k�$�2�������F�N��U���u�u�u�u�w�}�W���Y���Z�D�����g�1�"�!�w�}�W���
����^/��N��H����6�8�;�{�}�W���Y���F�N��U���u�u�u�u�w�p����
����WN��
�����_�u�u�u��>����Y���F��T��:���y�u�u�u�w�}�W���Y���F�N��U���x�u� �u�>�3���Y����G	�N��Uʦ�6� ��!�4�}�Iϭ�����F��['�U���u�u�u�u�w�}�W���Y���F�N��ʦ�2�0�}�b�3�*����s���%��V��������u�z�+����Ӡ��P��D�����4�u�4��w�p��������u��C'�����u��6�;�#�3���Y����[	��h��'���4�!�4�6�$�)��������R��t�����6�<�0�0�6�}�W���Y����[	��h��1����9�1�!�"�W�W�������RF��X��<����0�3� �]�}�Z�������@"��V'�����4�0��!�]�}�Z�������@'��B��U���6�8�;�_�w�p����&�ƿ�P��x������6�8� ��1�}���T����X9��D/�� ���!�&�6� ��)�}�������V��C������4�!�0�6�-�����Ξ�OǻN�����<�u�4�u�]�}�W���?����z��V��H����6�;�!�9�8�G���T�ƥ�F��X�����u�%�'�u�6�}�}���Y�Ɵ�^��t��U���k��8�9��6�W���Y���F�N��U���u�u�u�u�w�}�Z����ƿ�W9��P��U���u�&�4�4�6�4�W���GӒ��VJ�N��U���u�u�u�u�w�}�W���Y���F�N��Xʼ�u�7�:�0�9�}�W���
����R��V��H����4�!�4�4�8����:����p��g��1���,�x�d�y�w�p��������RǻN��U���!��u�u�w�`�W�������|��N��U���u�u�u�u�w�}�W���Y���F���U���;�1�d�u�8�3��ԜY���@%��Q��U���u�k�&�:�1�����Y���F�N��U���u�u�u�u�w�}�W��Y���@��R
��Gʱ�"�!�u�u�w�}��������F�
P��4���8�;�y�u�w�}�W���Y���F�N��U���u�u�u�x�>�}����������Y�����u�u��6�:�(�W���D�ƿ�P��x��Y���u�u�u�u�w�}�W���Y���F�N��X��� �u�<�;�3�i�W������F�N������!�6�u�i�.����6����_7�N��U���u�u�u�u�w�}�W���Y���F��CN�����}�b�1�"�#�}�}���TӲ��
��CN������9��9�.�*����
������R�����:�'�&�:�3�3�W�������_�������x�!�<�2�%�)�Ͻ�����G�������'�2�!�4�8�3�W�������Z��Y��U���&�u�:�3�>�4����Y���[����ʶ�;� �0�u�9�)�ϓ�:�ƭ�WF��RN�����9�!�1�'�$�1�W���������C��U���u��6�8�"�}����ӕ��]��d����� ��!�4�>�}�Jϭ�����R
��R��]���4�!�4�6�2�<�P�������]��c"�