-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����A��s������9�{�=�]�p�6�������\��v�����_�x��<�>�<�W�������6��R1�A߇�x�u�4�0�w�l�=���Y����9K��C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�w�>�W��Hӥ��J��_�����;�9��&�%�0����:����A��X חXʔ�9��2�!�w�8�������}��X ��U���!� �0�!�w�3����ӯ��\��C�����x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�Z��Y����\��N�����<�0�6�9�"�<�����Ơ�]�������9�!�1�6�2�;������ƴF�N��U���3�'�0�6�w��Y���Y���F�NחX���u�u�u�u�w�}�4�������]��Y�����'�<�0�u�?�>�W�������V����U���1�7�u�=�$�W�Z���Y���F��Y�����u��9�1�!�1��������U��^����_�x�x�u�w�}�W���Y����f��[�����<�u�&�0�#�9�W���Ӓ����R�����0�:�,�<�w�.�ϸ����F�N��U���=�u�:�3�>�4�����ƨ�_��[��X���u��u�!�>�}����UӒ��]F��RN���߇x�u�u�u�w�}��������]��R��ʼ�u�&�1�_�z�p�W���Y���F��^�����0�6�9� �6�8�W����Ư�V ��T�����#�'�u�9�4�}����W���F�N��U���:�0�!�0�2�4�W�������Z��CN�����;�u�0�4�w�3����Y����_�CחX���u�u�u�u��8��������]��V�����1�<�u�1�%�.���� Ӓ����C��D�߇x�u�u�u�w�}��������Z��X��%���0�;�u�=�w�n��������Z��Y��ʧ�4�u� �u�z�}�W���Y���\ ��R��ʴ�u�0�9�4�w�5�W������V
�������;�-�u�:�1�4����W��ƴF�N��U����0�d�u�%�>����ӄ��@F�������;�4�0�8�;�4����Y����[�N���߇x�u�u�u�w�}����Ӈ����YN�����!�u�=�u�%�:��������Z��Y��ʶ�9� �4�0�]�p�W���Y����������<�!�'�:�6�8�W�������V��=C�X���u�u�u�u�w�5�W�����������U���1�<�u�=�w�4��������C	��C��U���u�:�0�<�w�p�W���Y���F��RN��%���u�:�%�;�9�s�W���
Ӆ��C	��Y��ʼ�3�'�0�{�w�}�W���Y���9K�N��U���u��0�%�'�1��������G��B	�����u�:� �0�>�}�W������KǶC�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�_�9�5�<�Ϸ�����\��=N�����0�0�&�1�;�:���O�ȭ�_]ǻ��U���0�;�8�'�4�.�������F��@��[���� �<�<�>�.������ƹ����ą�2�'�6�<�9�1��������R
��=N�����:�>��2�%�>�3�������P��C����u�u�_�;�>�$�1�������\��t��U���_�u�0�0�>�u�W�������U+��~ �����u�u�;�0�2�t�}������F�V<�����u�o�<�u�8�1���Y����R��R-��U���;�&�1�9�0�>�}���Y����r
��X��U���;�7�:�0�9�W�W���)����z��� ���2�0�}��:�<����
����@K��S�����|�u�x�u�e�s�E���Yӕ��V ��B��U���u�<�;�1�e�}�������F�N��F���_�;�u�'�4���������P]ǑV�����!�'�u��w�;�1�������\��t��U���u�u�u�&�0�<�W�������	F��v#�*���h��!�:�1���������p	��Q#��<���4�6�|�_�w�4����
����V��NN�7���f�
�u�h��)��������R��E�����3��8�;�#�3���s�ƿ�T��������0�3�<�2�}�W�������	[��V��N���&�2�4�u��8��������C��N�����;�o�u�4�$�f�W�ԜY����R
��z����� �u�u�!��2��������U��S�����|�_�u�<�9�1����=����F��G��U���
�:�<�
�2�)���Y����G	�UךU���&�2�4�u��)��������\��C
�����
�0�!�'�d�}�������9F��^	��ʦ�9��8�4�6�(�'���Y�ƿ�W9��P�����:�}�`�1� �)�W���s����Z��[N�����<�<�;�u�w�4����K�ƨ�D��^��O���:�=�'�u�i�z�P��T�Ɵ� H�=N�����9�&�:�3��1���
����WN��
�����e�u�h�}�#�8���Y���F�=�[��_�u�<�;�;�.��������Z��T�����1�g�u�:�9�2�G���D�Σ�[��S�R��n�x�u�g�y�h�Wϭ�����@'��t�����!�u�u�<�9�9�F�������V�S�����'�u�k�r�p�f�Z���H���l�=N�����9�&�=�&�����Cӕ��]��\ ��6����4�0�<�$�l�W������F��F�����u�k�r�r�l�p�W��W���@��V��%���0�;�<�0�w�}����ۍ��^%��T>�����!�x�g�1� �)�W���C����G��DN��U��|�u�x��e�l�Wϭ�����@6��D��%���g�o�&�2�2�u�9�������R��^��D���:�;�:�e�w�`�_������F�G�X���d�{�_�u�>�3�ϭ�����]6��R]��U���;�1�>� ��1�'�������W��S�����|�o�u�:�?�/�W���^���K�d_�D���u�u�_�u�>�3�ϭ�����V
��g��E��&�2�0�}�e�9� ���Y���F��C����u�e�|�u�z��D��H����Z��[N������9�4�<�2�}�W������F��@ ��U���o�u�:�=�%�}�I���^���F��@��D���u�u�_�u�>�3�ϭ�����P��C>�����u�<�;�1�e�}�������	[�X�����k�r�r�n�z�}�E��L����Z��[N�����<�<�;��'�l�Mϭ�����T��X����u�h�}�!�2�.�J���I����K��]�@���&�2�4�u��8��������C��N�����}�g�1�"�#�}�^��Yۉ��V��
P��E���u�x��f�z�W�W���
����_F��B��Oʦ�2�0�}��:�<����
����@M��S�����|�o�u�:�?�/�W���^���F�=�[��_�u�<�;�;�.����Y����V��y�����=�&��!�|�}�������	[�X�����k�r�r�n�w�p�$��T���FǻC�0���'�u�=�!�#�8����8����V ��^��U���;�9�u�'�w�2�W���������XN��ʦ�2�4�_�u�z�����Y�����������0�&�4�0�w�8��������U����U���u�9�6�u�%�}����Y���\��Z��ʼ�!�u��f�$�}����������GN����;�n�u�4�#�4��������\ ��b�����0�3�<�0�m�.����Y���G��UךU���'�7�!�u�2�-����,����G%��Q�����u�<�;�9�>�}����[���R��^��ʾ�0�u�3�&�?�.�>���	����@��V�����'�0�n�u�6�)����Ӎ��CF�������0�!��%�g�}����ӏ����RL�Uʴ�!�<� �0�<�8�W���
����U��R �����o�&�2�4�w�.�U�����ƹ��E�����0�%�:�u��8����Cӕ��]��^�����w�_�u�u�z�+����
����R��N����>�&�2�;�]�?����s���6��R��ʴ�1�'�%�<�6�8����8����V ��C�����0�3�;�:�#�}��������R��R-��\���7�2�;�u�w�4�W�������W��d�����>�u�=�;�w�}�Wϭ�
����p	��Q>�����h�&�&��#�2���Y�����R/��6���3�<�0�u�j�.��������U]ǻN�����3�_�u�;�w�/����B���K��Y��U���u�:�3�<�>�3�W������ P��UGךU���6�&�}�4�'�8����Yӄ��ZǻN��ʧ�&�;�
�1�2�����:���G��N��U���u�x�u��6�8�Ϸ�Y����_F����U���4�0�6� �w�}�;���
����U ��S�����<���u�w�}�Z���)����z��DN�����u�:�0�u�?�3�F��UӒ��A��E��ʺ�9�u�0�1�#�8�F�ԜY���K��R��U���;�3�6�;�w�3����Y����FǻN��U���8�4�4� �w�`��������\9��C��¦�=�&��}��0��������Z��N�����u��8�4�4�5��������O�=N��U����8�4�4�"�����Dӕ��^"��V!��N���u�0�1�<�l�}����	����@��N�����x��0�3�4�8�Ϸ�Y����AF�������0�!�u�:�9�%�W�������V��^�����u�f�7�!�]�}�4�������]������&�0��!��)����J�ƨ�D��_�\���_�u��0�1�8����Dӕ��]��D#��1����!�<�0�f�}�������FǻN��U���x�u�;�0�w�5�W�������VF��R�����!�8�8�'�w�n�W���s�Ƽ�\��DF������>�_�u�2�4�}���Y����Z��P1�����4�%�0�9�~�)��ԜY���@'��z����� �u�h�&�;�����Q����]��R��%���0�;�>� ��1�'�������U��X��ʾ� ��9��6�8����H���l�N������8�4�4�"�����Dӕ��G+��s��:���_�u�u�;�w�;�}����Ƽ�\��DUךU���u�u�x�u�8�;�����ƥ���R��Fʷ�!�y��9�6�)�W���Ӆ��U ��^��U���9�"�'�d�w�4����
����\��^����u�<�;�1�$�1�:�������G6��RF�U���;�:�d�|�l�}�Wϭ�����U ��[��I���<�;�1�&�;���������Z��\�����:�e�|�u�w�W�W�������`��[���ߊu�0�<�_�w�}�Ϭ�
����V��=�����9�|�!�0�]�}�W���TӶ��V
��RN��ʳ�4�!�:�4�w�<�ϱ�Y����@��g��U���!�4�u�!�;�3�ϫ�Y�����������:�1�;�_�w�}�W������F��C�����!�<�u�0�3�}�ϼ�Y�ƿ�T���� ���;�:�1�'�#�}����Y����w5��+�����6�9�_�u�w�}�'�������C��S�����1�r�r�s�$�5����Q����p��g�����&�d�u�:�9�2�G���Y���F�D>������%�d�i�w���������]ǻN��U���4�0�;�<�2�}�Jϭ�����]6��R_�U���u�x�u�=�8�8��������[��V�����3�6�0�!�3�1�Ͽ�Ӓ����R�����:�3�<�<�9�}����s���F�:��ʥ�%�9�;�u�#�:�W���ӄ��[����U���<�2�7�!�2�3����;����R��C��1���m�u�9�6�]�}�W���ە��V'��t�����0�|�!�0�]�}�W���Y����U ��[�����u�h�&�9��8�������9F�N�����u�u�u�u�$�2��������C��S��6���3�0�!�n�w�}�W�������U]ǻN��U����:�&�u�2�*�����ơ�Z��X�����;�u�;�u�?�}��������P	��Q�����u�u�u�x�w�4����Ӓ��%��Q�����u�;�u�-�%�}����Y����VF�������4�0�3�'�#�8����Ӌ��G��^�����,�u�u�u�>�u�"�������U ��G��U���;�u�u�u�w�.��������G6��R^��Hʦ�9��0�3�4�8����Y�����Rd��U���u�&�:�3�>�4����	���F��X�����;�n�u�u�w�}������ƹF������6�0�!�<�2�}�J���:����Z��Y����u�u�u�0�3�4�L�������A	��D�U�ߊu�x��0�1�1����Ӗ��P����ʼ�3�'�4���e�������z ��_�����<�u�:�<�>�9�������K��_��&���9�8�;�u�$�4����������E�����u�%�:�0�$�����:���F��P��U���<�u�<�<�0�8��������p
�������u�u�x�u�;�}�Ϫ�ӂ��RF��G��U���u�0�<�!�%�9�����Ƹ�VF��gZ��U���=�9�u�<�?�)����s���F��_��<���%�f�i�u��<��������FǻN��U���0�3�0�!��-�F��Y����U ��[�����n�u�u�u�w�.��������G6��R\��Hʦ�:�3�<�<�9����Y���F�N�����u�=�u� �#�-����Y����~��R�����3��9�4�>�8�W���)����z��G�U���u�g�{�d�]�}�W���Tӥ��R��C�����'�u��!�w�5�ϩ�Y������Y�����0�7�!�u�1�)�ϰ�����9F�N��4���i�u�0�<�2�.����
����_��C��^����0�3�6�2�)����Y�ƿ�T��������1�9�;�#�}�W�������Z��g��G͹�;�!�|�|�]�}�W���Y����F��SN�����&�_�u�u�z�}��������[��B��ʺ�0�8�'�u�>�8�Wϊ��Ƽ�C��Y�����u�&�=�'�w�2�����ƾ�F��Pd��X���0�4�u�0� �8�W���
Ӣ��^��U��ʴ�1�!�0����'���Y����Xl�G�����4�0�0�y��0�������Q��Yd��Uʼ�u��&�!�#�8�}���Y�ƿ�\��x��I���:�=�'�u�i�z�P��Y����_�������0�2�}�4�'�8��������F�N������!�i�u�>�3�ǭ��ο�W��^	�����!�u��1�?�:�Z��P���F��SN��N���0�1�%�:�2�.�}���Y���F�=��U���n�