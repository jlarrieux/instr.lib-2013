-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����A��s�����;�!�:�!�8�s��ԑTӧ��[	��$��ʔ�8�'�4�_�z������Ɯ�\��CT��-���`�a��x�w�<����Oӫ��T��d����x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�Z���P����F��G������!�:�4�w�3��������p	��X�����x�u�9�u�>�5�ό�
����Wl� �����9��&�'�:�3�ϗ�����_F��Q�����;�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���6��G��O���=�&�3�9�w�0��������[��X �����;�!�3�'�#�8��������_F��T�����x�u�u�u�w�}�W�������]��Y��Uʐ�6�u�'�6�$�4�ϫ��ƻ�_
��V�����:�;�6�;�%�1�}��Y���F������u�=�u�:�#�2�W����Ƹ�_
��C�����u�3�!�0�'�2�����ƹ�Z��_�����u�u�u�u�w�<��������\��R��U���7�u�!�'�{�5� ϳ��Ư�P
����U���6�9�!�:�w�p�W���Y���F��[�����;�0�u�;�w�5�Ͻ�����Z�������4�0� �0�w�2�W���Y���F�N��Uʶ�9� �4�<�9�}�>�������R
��[��ʡ�0�&�4�!�'�<�ϸ�Ӓ����CNחX���u�u�u�u�4�3��������R��C��ʼ�u�=�;�!�w�)�����Ƣ�K��V�����:�{�x�_�z�}�W���Y����@��e�����!�u�:�6�w�5�W�������F�������'�u�=�u�"�/��ԑT���F�N�����9�!�:�u�9�}�����ƪ�AF��Y�����u�u�u�u�w�}�Z���Y���F�d�U���u�u�u�u��<��������GF��[�����6�;�'�9�5�2�϶�Ӌ��[F�������;�u�=�u�z�}�W���Y���P��R �����0�6�u�0�w�<��������9K��C��U���u�u�u�� �.�4�������K ��c��8���u�&�&�7�%�>��������[��B�����=�&�_�x�w�}�W���Yӄ��\��U��ʦ�;�u�=�u�%�>�3�������R
��N�����&�1�;�u�8�)�������F�N��U���:�3�<�<�9�}�����ƥ��������!�4�1�0�$�'����Ӓ����X�����x�u�u�u�w�}�W�������p	��Q'�����'�=�&��w�8�����Ư�]��[N�����3�!�0�6�%�8���Y���F�N�����6�0�!�&�8�1�W���
����P��U�������:�u�2�)�����Ƣ�K�CחX���u�u�u�u�$�<��������]��Y�����u�=�&�7�8�6��������P��R��ʦ�:�9�u�%�9�W�Z���Y���F��V�����;�u�0�:�2�4�W����Ƹ�VF��V�����=�u�0�!���Wϗ�Y����9K�N��U���u���=�$�;�����ƭ�_F����U���3�<�<�;�$�u����
�Ƹ�VF��E�����u�u�u�u�w�}����Y����A��R�����&�<�=�&��8��������g��z/��U���;�!�<�u��W�Z���Y���F��^�����9� �!�9�#�4�W���Y����P	��[��ʴ�9�:�u�!�w�<��������K�N��U���u�,�9�&�]�p�Z���Y���F�c�����9�;�u�0�6�}����
����G6��D�����!�u��-��>����6����_��C��U���u�u�u�&�2�(�Ϫ�Y����P%��[������0�~�d�]�p�Z���Y���F�c�����9�;�u�0�6�}����
����G6��D�����!�u��&�6�)�������K�N��U���u��9��6�8��������@F��T��ʶ�6�0�{�x�]�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���l��^�����0�0�u�:�<�W�W���Y������h�����d�a�4�9�]�}��������F��^�����9�n�u� �2�4��������P9��S@���ߊu�&�u�:�<���������Z��D����u� �0�"�%�s��������]��R�����{�9�n�u�]�3����?����w��E�����:�!�:�u�$�W�W������F��R��U���o�<�u�:�;�<�L���Yӵ��C
��[��U���&�1�9�2�4�W�W���Y����a��V��U���u�;�7�:�2�3�}���Y�����V�����8�;�u�u�9�(�����Χ�F��V�����d�1�"�!�w�t�W��,���l�N�����!�:�3��3�%��������\��YN�����0�}�d�1� �)�W���Y����T�d��Uʦ�<�=�&��2�;����?����Z��tN����;�<�;�1�f�}�������F�b_�D�ߊu�u��9��>��������VF��^ �����;�1�b�1� �)�W���Y����H��N�����u��4�!�?�.�!�������]F��X���ߊu�u��4�#�5����Y����]��Y������4�0�<�$�l��������F�;�[��u�u�_�u�w���������V)��a����:�!�7�:�2�3�}���Y����G+��g�����u�u� �u�9�4��������[��u��X���:�;�:�e�l�}�Z��W��ƹF�N�����!�'��9�w�}��������]]ǻN��6����4�0� ��1�������\	��V �U���&�4�6�=�$��������]��Y������9��4�2�4�������\F��U��Xǀ�f�d�_�;�w�/��������f��t�����_�4�6�<�2�)����-�ƣ� ��T�����6�;�!�:�#�2�W���Y���K��X�����0�u�3�!�2�.����
����_F��RN�����1�!�u�0�"�8��������F��YN�����<�0�_�u�>�3�ϭ����$��[��#���:�}�u�:�9�2�G���D�Σ�[��S����|�u�u�_�w�4����
����R��^��Oʷ�:�0�;�o�w�/��ԜY����Z��[N�����,�9�&�:�9�}�W�������Q��X����u�h�}�!�2�.�J���I����K��@�Uʦ�2�4�u��6�8����Y�ƹ�@��R
��;���=�&��!�z�}�������	[�X�����k�r�r�n�w�p�E���K���F��P ��U���-��6�=�$�����Cӓ��Z��SF�� ���4�0�<�&�f�9� ���Y���F��C����u�e�|�u�z��D��s�ƿ�T�������6�=�&��#�3�Mϼ�����l�D������-��6�?�.�8�������\��X����_�u�u�u�$�:����:����[��x������8�u�u�8�1����DӀ��@��N�����u��&�4�#�<����	����\	��V ��Hʳ�9�0�_�u�>�3�ϭ�����P6��D�����<��9�o�5�2����C�ƪ�_��=N�����9�&�0�!�%���������\	��V ��Hʳ�9�0�_�u�>�3�ϭ�����R��B�����6�u�u�:�;�<�W������l�D������9��4�2�(�;���Cӓ��Z��SF�� ���9��4�0�>�.�FϺ�����O�
N�����&�h�u�e�~�}�Z�J����Fǻ�����&�0�!�'��1�;��������[��U��3�9�0�_�w�4����
����c��R!��#���1�6��%�w�}�������� ��D�Uʦ�2�4�u��;���������c/��T�����;�1�>� ��1�'�������W��X����u�h�}�!�2�.�J���I����K��]�G���_�u�<�;�;�.���� ����~��D!��%���u�u�;�<�9�9�@Ϻ�����O��C��[�ߊu�<�;�9�$�<����	����\��X����u�_�u�!�%�?���������^ �����x��&�'�w�5�Ϫ�����Z��[N��U���u�0�2�1� �)�W�������A	��X��ʅ�'� �<�&�$�}������ƹK�E�����1�9�,�<�w�5��ԜY����Z��RN�����3�&�0�!�%����
����_F��L�� ���_�u�u�u�w�}�Z�������F��C��U���u�;�<�<�"�1����ӕ��]����U���u�%�<�<�2�}��������Z��[@ךU����<�u�<�;�5��������R��B�����2�<�&�0�y�}����������GN��U���9�o�&�2�6�}�������9F��C�����u�0�%�:�w���������Z��x �����u�<�;�9�>�}����[���FǻC�����
�<�&�4�#�}�Z¨�����Z��Sd�����_�u�%�:�2�.�����ʟ�^��t��U���7�2�;�u�]�}�W�������GO��_��U���u�&�1�0�k�}���������RG�U���u�&�0�!�%�����DӒ��V]ǻN��U���9��6�0��(���YӒ��F��P ��]����9��6�2���������[O��N��Uʦ�=�&��6�:�a�WǱ�����X�I����u�u��-��>����8����Z������h�u�e�|�]�}�W���7����R��V�� ���u�h�!� �l�}�W���
����~��_��:���;�<�0�i�w�/��ԜY���@(��C#��%���0� �u�h��)����D���O��N��Uʦ�4�6�=�&��)����-����[��V��N���u�u�&�0�#�<�'�������R
��{��I���4�&�n�u�w�}��������R
��R��I���4�&�n�u�w�}��������R
��T��Hʳ�9�0�_�u�w�}�4���)����|��V��9���i�u�4�&�l�}�W���
����c��R!��9���i�u�:�=�%�}�I���^��ƹF������!�4�6�6��-�W������l�N�����6�=�&��#�<��������Z�Q���ߊu�u�u��;���������c��R��]���0�&�h�u�g�t�}���Y�ƿ�R
��N����� ��0�<�2�a�WǱ�����X�I����u�u��9��0����Y����R
��dךU���9�<�u�<�>�:����Q����_��\G�����u�u�u�x�w�4����ӕ��@��CN��U���u�:�!�;�y�}�W���
����R��^��I����&�4�!�]�}�W����ƿ�V��E�����=�;�u�u�w�}�������	��R��H���'�0�n�u�w�}������ƹF������6�0��;�$�3�'���Y����p��t�����;�&�;�n�w�}�Wϭ�����^��C��Hʦ�4�6�,�9�$�2����Y����P%��[������0�<�0�]�}�W���TӢ��R�������0�!�_�u�w�}�9���4����R��B�����6�u�h�3�;�8�}���Y�ƿ�V��E�����8�u�h�3�;�8�}���Y�ƿ�R
��_��:���4�<��8�w�`������ƹF�C�6��� �4�0�!�2�?����Ӆ��G�������u�&�;�u��1�_���Y�����D'����|�!�0�_�w�}�W���TӢ��D��V��ʣ�9�1�&�4�#�-����Yӯ��@	�D��ʴ�6�9� �4�>�3�}���Y���K��QN�����'��%�u�$�<�����ƥ�]	����U���4�!�=�&��1��ԜY���F�������=�&��9�3�<�ϰ�ӕ��@��C>�����=�;�u�u�w�}�Wϭ�����G%��T:����u�'�0�_�w�}�W���Y����P6��D�����<��8�u�j�)���Y���F������h�}�!�0�$�`�W���
����F�N�����<�n�u�u�w�}�Z���Ӈ����C�����0�&�;�u�#�)�}���Y�Ʃ�@�N��U���u�u�u�&�6�>����6����_��R��I���'�0�_�u�w�}�W��8����VF��Y�����!�0�6�9�"�<��������@l�N��Uʼ�}��9��:�1��������F�N��Uʦ�1�0�i�u�8�5����GӒ��VO��N��U���u�&�0�!�6���������Z��[N�U���0�_�u�u�w�}�������F�R ����_�u�u�u�z�}��������@%��T-�����:�;�u�&�9�}�>���Q��ƹF������0�d�|�!�2�W�W���Y�ƿ�R
��N�����;�u�h�!��3��������p��t����� �!�9�;�#�t�}���Y�Ʃ�@�=N��U���u��9��4�8�4������@%��T-�����:�;�u�u�l�}�W�������U]ǑN��U���u�4�6�9�#�}�'�������^F��^ �����0�g�_�u�w�}�ǭ����O��_��U���u�u�&�=�$�����E�ƿ�G��g���ߊu�u�u�9�2�}�W���Yӕ��R��T��U��&�=�&��4�0�\ϭ�����]��Z��N���u�u�0�1�>�f�}���Y���%��T������-��6�?�.�6���ӓ��]��~
��]���u�u�u�x�w�2��������D��Y�����0�&�0�!�6���������G	��d�����&�u�u�g�}�.����0����^��@��U���&�u�u�u�z�}�Ϻ��Ʈ�P��RN��U���0�<�0�&�2�)��������P��X �����u�<�0�7�1�/�W����ƿ�]��XN��ʻ�-�u��{�w�}�W��Y����G+��g����� �u�&�4� �$�W�������	�������=�4�u�3� �8�Ϸ�Y����_��RN��U���:�8�1�!�w�5����Y���F��C�����9�;�u�!�0�s�W���Yӏ��@/��RF�\ʡ�0�_�u�u�w�}�9���4����R��T��U��&�!�'��6�8�\���)����z��R��¦�=�&��6�2�8�ȶ�����W	��C��\��r�r�n�u�w�}����s���F�D ������4�0�6�"�}�Jϭ�����P6��D�����~�&�=�&��>�������F�R ����_�u�u�u�z���������[��C�����u��r�u�?�.�W���Y����_��RN�����1�u��;�2�.��������@��C+�����0�<�!�'�3�W�W���Y����}��z������!�"�9�w�)�ϫ�����TF��T��ʼ�u�'�4�0�w�5�ϭ�����G%��Q�����:��<���W�W���Y����G+��g������u�h�&�2�)��������P��\ ��%���0�<�&�d�3�*����7����R��^�����=�&��0�1�3��������~'��[�����i�u��2�2�)����0����u	��_��4��_�u�u�u�z�����Y����U��[N�����4��4�0�"�W�W���Y����}��z������!�;�u�?�3�W���Y����}��z������!�i�u��%�:�������P��d��U���0�1�<�n�]�}�W���TӶ��V
��RN�����4��4�0�"��W���Y������Rd��U���&�0�!�4��<����<����VF������6�=�&��#�3�}���Y���F��G�����0�!�'��;�}��������R��B�����4�4�;�!�w�2��������\��_�����u�<�0�<�2�.�����Ə�_��V�� ���0�:�{�u�w�}�Z�������R��B�����&�:�9�u�$�8�Ͽ� Ӓ��VF��R�����9��9�4�$�/����0�ƿ�\����ʴ�&�'�u�;�#�0�W�������@��C8�����8�_�u�u�w�p��������]��RN�����:�0�6�0�1�>����Y����R
��[��U���=�!�<�u�8�)�������p��g��ʼ�u�0�&�!�6�}�ϻ�����\l�N��X����2�0�!�8�;�>�������[��v-��Uʜ�u� �;�u�"�}��������P��U�����8�;�1�7�w�����
����c��R!��#���1�0�u�<�?�}�W���T�ƿ�V��V����� ��u�'�$�8����)����|��Y>��ʦ�;�0�&�0�#�<�'�������^F�������3�&�=�&��>�ϼ�Y����P
��\N�����{�u�u�u�$�8����:����P
�
N�����'��9��:�f�W���Y����p��g������9�1�6�w�`��������R
��R�����&�4�6�=�$���������CF��SN��;����6�=�&��)�ϱ�Y����G+��g�������%�|�l�}�W���s���F�>�����0��9��6�8��������R��D�����u��"�&��8��������g��z/�����_�u�u�u�z�4�Ϩ�����\F��V�����6�;�'�9�w�3�ȭ�����Z��Y�����%�6�;�&�6�)�������F�N�U���u�<�0�<�2�.����Y������G�����!�8�;�u�.�.��������[��V�����:�u�3�_�w�}�W��
����c��R!��U���:�!�:�%�%�.�}���Y�ƿ�R
��_��:���6�u�h�&�?�.�6������F�D-�����&��!�6��-�W��
����c��R!��9���>� ��4�2�4�������\F��B�����<�&�&�4�4�5��������_��C��X����"�&��2�;����?����Z��tN�� ���2�0�}�0�8�u�4���)����|��T�����=�&�:�0�#�2��������A2��D#��R���2�=�|�n�w�}�W��Y����JF��RN�����3�!�0�:�#�(�ϱ�Ӆ��_��XN�����!�0�%�%�;�3�W����ƥ�9F�N��Xʴ�4�9�=�&��)����	��ƹF������!�4�6�6��-�W��
����R��V����u�u�u�u�$�<����
����e��S"��%���u�h�&�4�4�5��������W*��d��Uʰ�1�<�n�u�2�9��������9F�N�����u�=�u� �'�)�}���7����R��V�� ���9�1�i�u��%�:�������F��[����u�&�0�!�%�����Dӕ��@��C-������%�n�u�$�<����
����e��SN�U���9��4�0�"���������V]ǻ�����4�0� �u�j�.��������F��[>���ߠ0�1���]