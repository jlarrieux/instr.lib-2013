-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����A��~ �����:��:�>�8��!������r��X�?���u�8�0�8�9�p�W�������6��]��Oʅ��
�c�`�]�p�3���C����y��\�D���_�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z�ԑT�ί�T��N�����2�!��!�8�<�W�������]��t�����<�;�x�u�;�}����
Ӵ��V��Sd�U���<�;�9��$�/����
ӯ��V��[N�����4�<�;�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T��ƴl�>�����o��<�u�>�8�����Ƹ�R��V��U���8�!�0�&�3�1����	������CN�����u�u�u�u�w��W�������Z	��y��U��� �'�1�!�w�5�W���T����_	��TN�����:�u�=�_�z�}�W���Y�Ɗ�R��Y�����6�9�6��'�W�Z��Y���F�=��ʦ�2�4�&�4�2�4����ӏ��G��N��6ʶ�&�{��0�>�-��������QǶN��U���u�u�&�1�6�9��������G��^�����:�;�6�0�w�2�Ͻ�����GF��:��ʦ�8�_�x�u�w�}�W�������@F��RN�����u�;�:�4�%�$�W������5�����߇x�x�_�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���KǑ[�����<�0�y�"�%�f�Wϫ�ӏ��VH��S1�����d�c�{�9�l�}��������]��E�����4�9�_�u�$�}����)����f��^�����{�9�n�u�"�8� ���W����A��~ �����9�n�u� �2�*����������dװ���!�u�'�6��)��������P��G=��U���u�2�;�'�4�W�W���*����V��E-�����u�;�<�!�0�/�M���B�����R�����4�!�'�o�>�}��������U�=N�����_�u�u���:�%�������]F��S1�����_�u�u�4�'�8����Y����G��X	��N���u��0��<�g��������T��=N��U���0��&�!�m�4�W���&����P]ǑN�����6�;�7�0�9�g��������T��=N��U���!��4��3�8����
����\��YN�����2�6�#�6�8�u�W������]�N��[�ߊu�u��!��<�6�������U��N��U���&�1�9�2�4�+����Q�ƨ�D��^�U��� �{�_�u�w����������D�����6�#�6�:��e��������F�=�[�ߊu�u��4�2�3�W���ƿ�W9��P�����:�}�m�1� �)�W���Y����_�=d��Uʦ�4�4�;�4�>�}�W���
����\��d��Uʦ�4�4�;�e�m�4�W���&����P9��T��]��1�"�!�u�~�}�Zύ�A��ƹF��s��<���u�u�;�&�3�1��������AN��
�����e�n�x�u�f�s�}���Y����R/��N����!�
�:�<��8����H�ƨ�D��^�U����m�d�u�w�.���������D�����6�#�6�:��j��������F�=�[�ߠu�u�&�6�"���������\��D�����6�_�u�u��>����0����\��D�����6�#�6�:��h��������F�N��C��u�u�&�6�"����CӉ����h�����0�!�'�a�w�2����I���K��X����u��6�8�"��W����ƿ�W9��P�����:�}�`�1� �)�W���Y���`R�� d��Uʦ�6� ��!�f�g����
����\��h�����a�u�:�;�8�m�^���T�Ɵ�H��R ��3���!�;�0�%�%�>����-����e]ǑV�����!�'�u��w�;�1�������A��X�����:���<�]�}�Z���������V��ʡ�u�4�>�!�2�0����*����]��D@�����'�4�u�<�2�4�}���Tӂ��V��Y�����=�u�4�<�"�}����Ӊ��`6��D�����1�:�u�=�w��9�ԜY����R
��s��4���,�;�u�u�>�3��������GN��S�����|�_�u�<�9�1��������J/��T�����1�m�'�4��u�W������]ǻ�����&�=�&��%�$���)����l�
�����e�n�u�&�0�<�W�������W'��E��:���0��u�u�w�3��������R��_�����:�e�n�u�$�:����8����|��d�����!��!�#�l��������l�D������6�8� ��4����Y����|��CF����!�u�|�_�w�4����
����^)��a�����9�u�:�9�6�f�}���T����X9��P���ߊu�x�=�:��4����s����]l�C�����!�0�8�9�>��4ύ�/ӏ��F��^ ��U���4�'�,�u�9�$��������9F�N�����0��'�,�;�}��������]F��RN�����"�9�u�0�4�3�������F��@ �����u�:�4�:�3�(����
���� ��d�����4�'�4���a�Wǭ�����@"��V'��D���<�;�1�&�6�<���P���@"��V/������i�u�&�0�8�_�������O��^	��¦�4�4�;�e�~�W�W�������A��YN�U �&�2�0�}��<����Pߓ��Z��SF������e�|�_�w���������A��x�����u�u�h�}�9�4����
����a��v
�����3�&�!�|�"�.����Q����R4��S/������3�0�e�~�W�W��Y����A����U���'�%�<�!�w�/��������\��X�U���u�=�&�2�9�/���������������u�9�-�7�;�)�W�������\��@�����:�u�4�=�w�p�W������K��X��ʓ�4�!�;�0�'�/��������9F������u���2��.�Ϫ�&����V��V"�����0�0�|�u�z�+����ӕ��V��D�����:�9�4�}��8�%������K��X��ʦ�4�6�;�7�2�)�(�������@%��T+�����;�_�u�x�?�2�(���)������V������}��8�;�.�������W��X����_�u�x�=�8��W�������W'��E��:���0��u��#���������| ��R��]���8�9�&�0��>���Hӂ��]��GךU���=�:�
�u��)�>�������\9��X��¦�4�4�;�4�>�t�W������l��s��<���&�4�4�'�6��>ǵ�����@6��t�����d�1�"�!�w�t�W������l��s��<���&�4�4�'�6��&ǵ�����@6��t�����d�1�"�!�w�t�W������l��v������9�1�&�4�(�8�������\	��N����>�4�&�6�"�����8����|��d������8�9�&�2�����T����\��XN����x�=�:�
�w���������r��Z!��$���;�1�>�4�'�8�'��� ����F��S�����|�u��4�#�3��������\��X��U���<�,�"�'�y�/��������A	��[��!���}��|�u�w�:����Ӌ��NǻN��U���8�9�&�0��>���Y����C
��g�����y�u�x�<�w�4�������l�N�����'�9�6��4�2�W�������P
��\(�����u�x�u�;�w�3����Y���9F���ʸ�%�}�u�u�w�<��������GF�N��U���u�h�u�:�5�2��������T��D��Y���u�u�u�u�w�}�W���Y���F�NךU���u�4�%�0�;�}�W���Y���F�S�&���9��>�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�x��6���u�u�u�u�w�}�W���Y����E��[�U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���
����a��CN��U���u�u�u�u�j�}����������R�����y�u�u�u�w�}�W���Y���F�N��U���_�u�u�u��1�2������F�N��U���k�!�
�:�;�<�_�������Q
��YG�U���u�u�u�u�w�}�W���Y���F�N��Uʦ�=�&�u�u�w�}�W���Y���F������'�4��}��0��������_�_�����:�e�y�u�w�}�W���Y�����C��#���1�u�u�u�w�}�W��Y����\	��V ��1�����9�1�{�}�W���Y���F�N��U���u�u�u�_�w�}�W�������W'��E��:���0��u�k�$�<��������V��Q�����>�4�%�0��/����Y����W	��C��\�ߊu�u�u��#��>���Y���F�N��U��&�4�4�'�6��>ǵ�����@6��t�����d�1�"�!�w�t�W���Y���l�N�����4�;�u�u�w�}�W���Y���X��s��4���,�;�}��:�1����:����K�
�����e�y�u�u�w�}�W���Y����r��Z!��#���1�u�u�u�w�}�J���8����|��V��7���y�u�u�u�w�}�W���Y���F�N��U���u�u�_�u�w�}�6�������F�N��U���u�u�k�&�4�(�8���*����WN��V�����'�,�9�u�w�}�������F�N��U���u�&�6� ��)�W���Y���F�N��U���6�8� ��>�3�ǵ�����@6��t�����d�1�"�!�w�t�L���Y��ƓF�v����� �%�!�_�w���������Z�S�����1�:�<�}��>����/����q	��UךU���6�8� ��w�a�W���&����P9��T��]���6�8� ��>�3���P���@'��B����u�h�&�1�;�:��������@'��B�����2�0�}�|�l�}��������zW�S�����:�<�
�0�#�/��������z5��Y��D���"�0�u��:�1����:����[������!�0�&�h�w�m�^�ԜY����F��C?�U��&�1�9�2�4�+����Q����F��C?�����}�|�u�=�9�6��������p��RN��Gʰ�&�u�:�=�%�}�I���^��ƓV��e:��