-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����A��~ �����:��:�>�8�s��ԑTӧ��[	��$��ʔ�8�'�4�u�9�}����:����]	ǶN�����4�u�'�?�4�g�'���&����al�*�����l��9�u�g�l�Z�ԑT���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���6�u�e�d��-����Ө��Z	��[N�����8�;�&��%�2�������r
��e�����0�0�#�1�z�}��������]��B�����;�0�;�9��;������ƴK�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���_�x�x�u�"�-���Y���� ��RN�����&�4�%�:�2�.��������U	��C�����!�:�4�_�z�}�W���Y����]��G�����u�!�!�>�$�4�W���Ӊ��G��d�����>�1�8�<�y�}���Y���F�N�����:�0�u�=�w�<�Ϫ�Y����|��t�����<�u�=�6�w�.��������WF��R���߇x�u�u�u�w�}��������p
��N��ʱ�2�!�9�&�0�<�W�������]��DN�����;�!�0��2����Y���F�N�����u�;�u�=�9�)�ϱ�����W�������&�0�'�1�5�>�W�������R��R-�����u�u�u�u�w�9����W���K�N��U���u��0�6�8�6����ӏ��Z��R�����4�,��0��6�����Ƹ�V��V��X���u�u�u�u�w�2�W���ӵ��C
��[�X�߇x�u�u�u�w�}��������C
��g�����u�;�<�4�2�5� ϳ��ƿ�^��DN�����;�<�,�x�w�}�W���Y�ƾ�P��R��ʡ�0�&�4�4�9�r�W������@"��V'��Z���'�u�4�&�3�p�W���Y���F��@ �����u�;�4�&�9�1�W���Y����F��T�����;�u�;�!�2�<�������F�N��U���4�&�1�:�w�}��������|��T��ʶ�6�0�u�:�w�5�Ϭ�����K�N��U���u��%�!�6�-��������VF��R
�����0�&�4�9�%�)����Ӄ��R
��Xd�U���u�u�u�u��8�4�������\�CחX���u�u�u�u��4�W�������G��DN�����6�9� �4�>�3���� Ӓ��VF��V�����0�x�u�u�w�}�W���
����@H�u��ʺ�u��4�0�w�)� ���Y������T�����=�u�<�!�%�2����s���F�N��U���6�8� ���2����Y������A��ʢ�0�u��6�:�(�!���Ӈ��V��N���߇x�u�u�u�w�}����Y����[��R
�����!�0�&�<�#�/��������JF��D�����&�4�4�;�6�4�}��Y���F���ʣ�9�1�1�!�w�4�W�������XF��T��U���0�u�;�&�6�<����WӲ����VחX���u�u�u�u�$�2����ӏ��_��Y��U���!�0��7��
�1���Y����A��=C�X���u�u�u�u�w�5�W����ƨ�G��R�����0�&�u�;�w�5��������[��
�����;�u�<�0�>�8�Z���Y���F�S��ʦ�'�6� �0�y�	�ϲ�����V��E�����;�<�0�"�.�)�W����ƭ�_F��Rd�U���u�u�u�u�6�5�[Ͽ�Ӂ����ZN��U���6�u�=�u��}����Y����[��V�����u�&�!�_�z�}�W���Y����V
���������<�u�?�}�!Ϛ�����F��V�����u�=� �1�%�<�Ϫ��ơ�W��=C�U���u�u�u�c��8�4�������@F��C�����6�;�7�0�w�3����ӑ��W��s��<����8�&�_�z�}�W���Y����VF��[����>�#�'�9�4�����Y����V��X�����u�=�u�0�#�2�W���Y����GǶN��U���u�u�<�u�?�}��������W	��^ �X���u�u�u�u�w�2�ϭ�����e��SN��ʦ�4�4�0�1�3�/��������]F��RN�����0�%�6�0�w�2�Z���Y���F�U�����4�<�;�1� �)�W�������_�u��U���!�<�u�<�9�1�W���Y����	��=C�U���u�u�u�6�4�8�����ƿ�R��Y'��U���u�!�<�u�8�}��������\F��A��U���'�9�_�x�w�}�W���YӅ��_��X�����u�;�!�0��}������ƴl�N��U���u�u�:�u��0��������_�\����4�0�1�1�%�.�8�������P	��V��U���<�!�2�'�z�}�W���Y���\ ��R�����!�u�2�:�2�)�ϸ�����R��R��ʡ�0�&�<�!�%�:����
�Ƙ�Z��Dd�U���u�u�u�u�2�9�ϼ�������*��ʶ�8�&�<�u�%�(�ϱ�Y����C
��g�����y�"�<�=�:�<���Y���F�N�����1�!�u�4�w�8�����Ƹ��������&�u�#�;� �8�W����Ƣ�GF��CN�����u�:�_�x�w�}�W���YӒ����E��U���6�9�!�:�y�����
����a��v
�����3�&�!�;�!�1�������D�^����u�u�u�u�w�<����I��ƴF�N��U���u�e�u�k��8��������GF��C�]���8�;�u�u�1�)�ϲ�
�ƺ�_��S��Y���u�u�u�u�w�}�W���Y�ƥ�P
��^ �����1�!�u�=�9�.��������WF��D�����x�u�u�u�w�}�W���H���f��C�����;�u�0�0�#�9���Q����V��N��U���u�4�!�#�;�9����U���F�N��U���u�u�u�<�4�(��������R��@��U���!���9�3�<����
��ƴF�N��U���u�d�u�k��8����������R�����{�x�u�u�w�}�W���Y���F��^��ʻ�!�4�#�9�3�2����W���K�N��U���u�=�u�:�"�8�����ƾ�@��@��U���u�&�;�=�8�2�Ͽ�����a��CN��U���4�&�'�<�0�p�W���Y���F��D�����{��<�u�8�(�Ϭ�����@F��D�����u�:�7�u�%�8����Ӈ��u��e�����u�u�u�u�w�}��������9K��C��U���u�u�u�=�w�4����ӂ��R��_�����=�&�8�1�;�}���Y���F�N�� ���%�}�u�u�g�v�F���6����_	��q�����~�d��8�;��Ͻ�����9K��C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�_�>�/�������D	��d�� ���<�0�{�!��2����H����_
��N��ʼ�0�{� �0�>�������ƹ����ą�2�<�!�9�#�8�3�������F��RN�����>��%�4�;�W�W���Y����6��q�����0�%�4�9�]�8����Y����G/��R�����9�6��%�>�W�W�������9F������&�0��6�2�g��������AF��_�U���>�#�'�9�4�����Y�ƥ���R	��U��f�n�u�%�%�u�W�������T��D��Oʼ�u�:�9�4�l�}�Wύ�����_������9�2�6�_�w�}��������Z��C
�����n�u�u�&�$�/����Y�ƥ���[��N�ߊu�u��9��<����Y����\	��V �U���&�=�&�u�m�4�W���
����X5��G��%���,�9�x�u�8�3���B���fT��dךU����!���;�9�MϷ�Y����V��=N��U���!��4��3�8����
����\��YN�����0�g�'�4��u�$�������A%��[��U���;�:�e�n�z�}�E��Y����w��~ ��Oʼ�u�<�;�1�o�/����Q����C
��g�����x�u�:�;�8�m�L��Y����l�N�����;�u�u�;��:���8����l��d�����0��6�0�f�9� ���Y����K��V����u�&�6� ��)����Y�ƣ�GF��X���ߊu�u��6�:�(�>������R��B��]���8�9�&�0��>�������\F��N�U��{�_�u�u��>����(����F��V�� ���}��8�9�$�8�4�������\��XN�\���x��c�b�2�9�1�������A��X�����:�n�_�'�?�)����Ӵ��	��q�����0�%�'�6�;�>�#�����ƹK�a��ʜ�!�'�:�4�>�3�1�������\��_�����9�u�'�u�w�3�W��6������B�����u�:�_�u�z�?��������l�D�������>�4�#�/����&�ƥ���R	��U���2�u�u�:�9�2�E�ԜY����V��NN�����9�6��6�8�}�Ϸ�Y����VF��Q��ʷ�u�#�9��4�2�%������F�:��ʴ�6�<�0�!�%�}����
����A��D��U���2�{�u�6�9�)����/����J)��[�����u�u�#�9��>��������9F�N��U���u�u�u�u�w�}�W���Y������R�����4�!�'�_�w�p�W����Ƃ�^����&���9�&��'��>�ϸ�Ӓ��@F��S��U���u�u�:�>�!�/����?����AH��C�����x�#�9�0�w�<�����ƻ�Z��YN��U���<�2�0���}��������[Hǻ�����u�%��;�2�)��������AF��Y	�����'�9�6��4�2�W������l�C�����,�>�4�%�2������ƥ���E��ʱ�3�;�1�7�w�-�%������F��Y������'�3��'�)����Yӵ��a��R1��U���u�u�u�u�w�}�W���Y���F��=��'���0�!�>�4�'�8�'��� ����lǻC�!���;�8�0�u�1�����
����f��DN�����u�0�6�%�5�8��������V��Y	ךU���>�:�,�=�$�����5����[F��[�����!�:�&�4�4�0��������V��N��[���x�u��8�%�>��������@F�t�����>�:�,�=�$�����5����[I��A������6�:�|�w�>�����Ƨ�F��X����� �<�&�o�9�)����Y���F�N��U���u�u�u�u�w�}�W��Yۍ��_��V�����'�0�2�=�|�6��������R��EN�D���u��0�6�8�6�������K��_�����=�:�u�=�w�2�����Ƹ�\F��T��ʢ�&�6�'�3�;�$��������9F�N������;�u�4�w���������P��E��U���u�;�u��#�(�$���Y����F������:�>�4�!�%���������V��[�����0�6�<�0�w�3����	����@ǻC����u�&�&�!�>�}������ƹ��Y�����4�;�,�6�m���������\��x�����>�4�!�'�3�*����P���	��R��H���4�&�|�_�w�4��������G5��TN�7���0�;�0�!�%�6��������R��EN�����u�|�o�u�8�5����GӀ��@�=N�����9�:� �%�#�$���;����R��T��]���0�6�:�>�6�)�������\F��T��]���0�&�h�u�6�.�^�ԶYӕ��]��D-�����7�0�<�0�m�?�������U��RUךU���;�9�&�4�6�3����)����	F��X����u�4�&�n�w�.����Y����@��G��U���&�
�}��:�1����:����W��X����u�h�}�!�2�.�I�������[�^��\���x� �l�m�w�.����Y����R4��S/������3�0���-�W�������V��E��*����8�9�&�2�����Hӂ��]��G��H���!�0�&�k��)����D���O�C� ���_�u�<�;�;�.��������zF��d�����'�,�!�<�<����)����P
��N�����u�|�o�u�8�5����G�Σ�[��S�E���n�x�u�d�y�W�W�������w��~ �����o��2�0�f�����ۍ��^��D>��6���0�d�1�"�#�}�^��Yۉ��V��
P�����'�u�k�e�~�f�Z���H����9l�D������9��4�;�}�W�������	[��V��N���&�2�4�u��)�>��������[��U��3�9�0�_�w�.����Y����R4��S/������3�0��w�}��������A��h��&���9�&�0��4�8�FϺ�����O�
N�����&�k�}�!�2�.�J���I���K�b\����<�;�9�:�?�.�W�������GN��V�����'�,�9�x�w�2����I����N��_��H���:�=�'�u�i�z�P���Y���� V�=N�����9�:�4�4�9�}�W�������r��N1�����%�0��'�.�1�Z�������V�S�����'�u�k�}�#�8���^���F�=�[�ߊu�<�;�9�8�<����Y�Ɵ�T��V�����!�>�4�%�2���������W	��C��\��u�:�=�'�w�c�_������A��G�X���d�{�_�u�>�3�ϱ�����`��V��Oʦ�2�0�}�b�3�*����P���	��R��H��r�n�x�u�f�s�}�������	��C��&���4��o�&�0�8�_������\F��T��]���0�&�h�r�p�f�Z���H����9F��^	��ʺ�!�'��9��)�Mϼ�����\�Q���ߊu�<�;�9�8�<��������R�������u�h�3�9�2�W�Wϭ�����\'��B�����<�o�7�:�2�3�M�������9l�D������6�8� ��1��������\	��V ��Hʳ�9�0�_�u�>�3�ϱ�����F��G��Oʑ�!��!�!�<�<����)����P
��N�����u�|�o�u�8�5����G�Σ�[��S�E���n�u�&�2�6�}�6�������Z��T����� �
�}��:�1����:����W��X����u�h�}�!�2�.�J�������@F�^��\�ߠu�&�2�4�w���������Z��[N����9�2�6�o�w�m�L���
����_F��T��:���6��o��#���������_��R�����d�1�"�!�w�t�M�������@F�F�����u�k�e�|�l�p�W��W���@��V��4���8� ��9�w�}��������X5��G��%���,�9�x�u�8�3���Y���\��E��K���!�0�&�h�p�z�^���Tӵ��QǑN�����u��!���9��������V��X	�����}��0�6�8�6����ڂ��]��G�Uʦ�2�4�u��9�����Y����T����G���&�}��0�4�2��������\��XN�N���&�2�4�u��<��������u\��X����_�u�4�!�>�(�ϳ�����\�������_�u�!�'�5�)�W���&����F��QN������;�u�u�>�3�Ϸ�Y���9l�C�����u�<�;�9�w�<�Ͽ�[����F��C�� ���!�u�;� �2�)��������\��	�����x�&�6�0�w�3�ύ�5�Կ�F��R�����&�!�u�0�6�3�W����Ƽ�G��R�����=�_�u�x��0����Ӈ��)��E-��U���4�;�u�:�w�4����s�ƭ�G��B�����u�u�!�<�0�W�W�������VF��R��ʺ�4�6�;�7�2�g�����ƥ�D��B�����!�'�7�!�w�8�ϱ�Y����R4��S/������3�0��w�}����ӏ����RL�Uʴ�!�<� �0�<�8�W�������z��[��Oʦ�2�4�u�&�u�/���YӇ��A��C�����:�u��4�2�g�����ƥ�D��B�����!�'�7�!�w�8�ϱ�Y����R/��T�����9�<�u�!�"��}�������F��\��U���:�4�4�;�w�}����ӏ����RL�Uʴ�!�<� �0�<�8�W���
����^)��a����&�2�4�u�$�����B����G��U��U���%�:�u��4�0����Cӕ��]��^�����w�_�u�!�%�?��������UF��T��:���u�u�<�;�;�4�Wͪ�����9F�N�����&�2�4�&�?�+�W���������E�����:�0�&�'�w�5�Ϫ��ƨ�]A��P��U���u� �>�1�>�)�W���J���2��E�����u�:�7�u�w�2����Ӗ��[F��C��ʡ�0�u�x�u�!�/�����Ɵ�^��t�����<�&�3�'�#�0���YӇ��A��C�����:�u��6�:�(�!���������Y�����!� �w�_�w�)�����Ƨ�V��QN������!�6��w�4��������A��d�����<� �0�>�2�}�ϭ�����F��[?����4�u�&�w�%�8�L�ԜY����]��RN�����=�u�,�6�'�-����Y����R
��XN��ʲ�!�<�%�0�2�)�ϩ��Ɵ���X�����2�u�4�!�>�(�ϵ��ƣ�	��G�����u�<�;�9�>�}����[���R��^��ʾ�0�u�3�:�6�<�����ƿ�T����W���0�n�u�4�#�4��������\ ��x�� ���;�o�&�2�6�}�������9l�C�����&�2�!�'�]�}����Ӊ��P��B��U���4� �
�}��0��������_�
�����e�n�u�&�0�<�W�������G7��s��:���!�>�4�%�2���������W	��C��\�ߊu�<�;�9�8�$��������Z��U�����_�u�x�=�8��������T��N�U���6�u�=�u�9�(�W�������Z��_�����0�9�u�:�6�3�����Ƹ�V��E�����!�_�u�x�#�8�8���:����\��Y@��!���u�&�1�;�w�2�����Ƹ�V��^��U���9�2�6�u�z�}��������V��_�����;�u�:�u�>�4��ԜY����V��V"�����0�0�y�4�'�8����Yӄ��ZǻN��´�#�%�4�0�2�t����s���F��V�����0�<�0�u�w�}�W������l�N�����4�;�4�<��-�W���Y��� ��D�U���u�&�=�&��-�W���Y���F�S�����'�h�u�:�?�/�W���^���l�N�����4�0�1�1�%�.�8�������Z��N��U���h�}�!�0�$�c�_������F�G����u�u��!������Y���F�R��]���0�&�k�:�?�/�W���^���l�N�����4�;�<�0�w�}�W���Y���N��_��H���!�0�&�h�w�m�^��Y����_�������0�2�}�4�'�8��������F�N�����;�7�0�<�2�}�W���Y����p��r ����u�u�u�&�6�<��������VF�N��I����!���;�9�}���Y�ƿ�R��R�����&��3�0������Y���Z�D*�����1�1�'�&��;����B���F��g�����0�u�u�u�w�}�W��Y����@��N��Uʦ�4�4�;�<�2�}�W���Y���[��s��<���_�u�u�u��)�>���	���F�N��U��&�4�4�;�l�}�Wϻ�ӏ��9F��Y
�����&�n�_�u�z���������]�������u�;�!�0��8�4�������]H�c��U���1�;�u�:�2�.��ԜY����[����ʻ�x�:�<�u�6�5��������[��X��ʳ�'�!�8�;�y�}����������P������0��>�]�}����s���Z ��{�����&�!�u�=�9�}�W�������v��[��Hʳ�9�0�_�u�w�}�3���0����Z�
N�����_�u�u�u��<���Yۉ��V��	N�����&�h�u�e�~�f�W���YӉ��G��V
�����&�3�&�!�9�a�WǱ�����F��C����u�e�|�n�w�}�Wϱ�����zF�F�����u�k�}�!�2�.�J���I���9F�N��1�����i�u�8�5����G�Σ�[��S�R��|�_�u�u�;�4�W�������W��x��6���u�=�;�u�w�}��������_�
N�����;�7�0�<�2�W�W���Y����R/��V��U��&�4�4�;�6�4�'���B���F��g����u��4�0�>�8�}���Y�ƣ�R��R�����&��3�0��}�Jϭ�����R��S�����&�!�;�<�2�W�W���Y����R/��R�����4�;�<�0�l�}�W�������z��S��1�����%��]�}�W���Y����F��SN�����&�_�u�x�w�/��������z��C=��ʦ�2�4�u�=�#�)��������E��[��3���=�;�!�u�6�-����T�ƨ�G��E������8�9��<�9����W�Ə�V����U���!� ��;�w�4��������G��Dd��X���=�u�#�'�;�}����Ӡ����YN��U���6�u�=�u�6�<��������[��B��ʆ�8�9��>�w�p�W�������u��R��ʶ�'�0�!�,�]�}�Z�������|��T������;�� �#�/�W������l��x�����>�4�!�'�<�+��������G	��N����>�2�>�:�9�������� V�N����>�4�4�0�2�}�;�������VǻC�����
�u�4�0�;�}��������F�A������0��>��8�4���Y����[	��h��6���!�:�,�6�8�3�}���T����X9��X-�����9�1�:�,�4�2������ƹK��_��*����&��>�3�8��������F��R�����;��;��"�)�������JF��E�����9�6�<�2�.�>��������g*�N�����'�6�8�%��}�W�������P
��\(�����h�u��0�4�2�������K�^ �����2�'�o�u�]�}�W���:����~��V �����k�w�e�|�w�}�W���Y���K��YN�����2�o�u�f�u�}�WϮ��ơ�CF�N��Uʴ�0�0�u�u�w�}�W���GӇ��u��e�����u�u�x�<�w�?�������F��V�����u�u�u�u�j�}��������F�N��X���;�u�!�
�8�4�}���Y�ƃ�V��\N��U���u�u�k��2�����Y���F�N��Uʦ�1�9�2�6�w�}�Wϱ�����F�N��U��u��;��"�)�W���Y���	�������1�9�2�9�$�l��������X ��C���ߊu�u�u��"�)����Y���[�X=�����;��9�1�w�p�W���Y����V��N��Uʺ�4�0�9��0�����GӉ��]O��N��U���u�u�x�:�#�?�������K��^�����!�0�&�;�w�4����Y����R��C�����4�<�'�!�w�8����0����`�������9�;�1�u�z�}�8�������u��X��U���,�9�&�u��)�����Ƨ�E��[��3���:�u�,�9�$�W�W��7����G���� ���<�u�:�u�.�>�Ϫ�Y����`��[��ʰ�2�u�8�0�>�)��������R*��G	�����{�u�x�u�?�/����Y����@��d��6���!�4�<�u�8�0�����ƹ�@��R
��6���!�6�8�4�>�2��ԜY����V��V"�����0�0�y�#�%�1�^�������9F������%�4�0�0�~�)��ԜY���\"��V'�����u�i�u�:�?�/�W�������]ǻN��U���%�!�,�6�w�}�J�������[�Q����u�u�u�:�"�-�������F��C����u�4�&�|�]�}�W���=����]/��R��I���:�=�'�u�i�z�P��Y����_�������0�2�}�#�%�1�^Ϫ����F�C�����0�9�u�;�"�}�����ƭ�VF��P�����u�<�&�u�9�)�ύ�����_��X�����u�u�x�u�9�}�����Ƹ�VF��R��ʱ�8�<�{��>�}����Y����p
��D�����"�9�u�0�]�}�W���TӒ��Z��R�����&�:�u�=�w�8��������\ ��A�����3�0�u�u�>�4����Y���F��P��ʆ�8�9��>�6�9����Y����AF��[�����'�9�6��4�2�W������F�N�U���u� �!�%�2��4Ͽ�Ӌ��V��Y��ʦ�;�9�u�<�9�1����Ӊ��]��B �����=�_�u�u�w�p����Ӈ��	��C��&���u�&�0�!�w�3��������@F��������8�9�&�2�����Y���K�^ ��U���u�4�4��:�/�Y���Y���F�������'�6�&�<�0�8����������RN�����;�0�"�u�6�6��������_��@�����u�u�x�:�9�(�$���s���F�:�����'�u�=�u�6�-����Y����Z��R�����u�4�<�u�"�-�ϸ��Ƹ�VF��T�����'�u�u�u�z�}�Ϲ��Ƹ�VF��C��U���;�9�u�&�9�}��������l�N��X�ߊu�u�u�x��/�W���ӂ��T�������&�'�!�u�8�}���� ����Z��[�����&�<�;�1�]�}�W���T���F�N��U���u�
�
�
��}�W���Y����l9��h1��U���u�u�u�
���(���Y���F��V�����u�u�
�)�w�}�W���&����l9��N��U���)�
�
�
��}�W���YӚ��l9��h1ךU���u�x�u�u�w�}�W���Y���l9�N��U���
�u�u�
�w�}�(���Yӹ��F��hN��U���u�u�
�u�w�}�Z���6����_�N��*���u�
�)�u��!�W����ư�l�K1��Uʩ�
�u�)�
�w�!�(�����ƹF�C�U���u�u�u�u�w�}�W���&����l9��h1��*���
�
�
�
���(���&����l9��h1��*���_�u�u�u�z�}�4�������WF��hךU���u�x�u�u�w�p�Wϱ� ����F��N��	���u�)�u�u�+�}�WϢ�Y����F����G���u�e�u�u�f�}�W��Y���F�C��U���u�u�u�u�w�}�W���Yӹ��l9�N��U���u�u�
�
�w�}�W���Y���l9��hd��U���x�u�:�;�"�����Pӹ��l9��KN��Uʩ�
�
�
�
��!�W�������l9��h1��U���u�
�
�
�w�}�W��Y���F�N��U���u�u�u�u�w�}�W���Y���F�h1��*���u�u�u�u�w��(���Y���K������,�6�=�2�~��(���&����l9��h1��*���u�u�u�
���(���&���F��h1�����u�u�x�u�w�}�W���Y���F��h1��*���
�
�
�
�w�}�W��Yӕ��_��V��Uʊ�)�u�u�u�w�}�W���YӚ��l9��h1��*���
�
�
�
���(���&����9F�N��X���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�
���(���&����l9ǻN��U���u��9��6�1�Wρ�&����l9��h1��*���
�
�
�
�w�}�W���Y���F�K1��*���
�
�_�u�w�}�Z���Y���F�N��U���u�u�u�u�w�}�W���Y���9��h1ךU���u�x�u��6�)��������l9��h1��*���
�
�
�
���W���Y����l9��h1��*���
�
�
�
�]�}�W���T���F�N��U���u�u�u�u���(���Y���F�1��*���u�u�u�u�w�}�(���s���F�N�����;�,�6�e�w�}�'���Y���O9��h1��*���)�u�u�)���(���&���F��h1��*���u�u�x�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���&����F�N��U���
�
�
�u�w�}�Z�������z��Y�����u�u��
���(���&����l�N��*���
�
�
�
�w�}�W���&��ƹF�C�U���u�x�u�u�w�}�W���Y���F�N��*���
�
�
�u�w�}�W���&����l9��N��Uʊ�
�
�
�
��}�W���T����w��~ �����|�g���+�}�W���Y����l9��h��U���u�u�u�
���}���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���
�
�
�
�w�}�W���&����l9��hd��U���x�u�:�4�6�3��������T��g-��*���
�
�
�
��!�W���Y�����h1�����u�u�x�u�w�}�Z���Y���F�N��U���
�
�
�
���(���s���F�N�����;�4�<�u��}�W���Y���F�N��*���
�
�
�
���(���&����l9��h1��*���u�u�x�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���&����l9��h1��*���u�u�u�x�w�2��������WF��h1��*���
�
�
�
���(������F�N��U���u�
�
�
���(���Y���l�N��X���:�4�4�;�6�4�0���s���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�
�
�_�w�}�W��Y���F�N�&���
�
�
�
���(���&����l9��N��	���
�
�
�
���(���&����F�N�U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�
���(���s���F�N��U���u�u�g����(���&����l9��h1��*���)�u�u�u�w�}����&����l9��h1��*���u�u�x�_�w�}�W��S���L�D��_�������}�w�]���S���L�D��_�������}�w�]���S���F�N�U���u�u�u�u�w�}�Wρ�&���F�N��U���
�
�u�u�w�}�W���Y����ll�N��X���:� �%�!�.�>�GƁ�Y���O9��h1��*���)�u�u�)���(���&���F��h1��*���
�
�u�u�w�p�W���Y���F�N��U���u�u�u�u�w��(���Y���F�N��*���u�u�u�u�w�}�(���&���F�N��:��� ��;�}�>�5�(���&����l�N��*���
�
�
�
�w�}�W���&����l9��Kd��U���x�u�u�u�w�}�W���Y���F�N��U���
�
�_�u�w�}�Z���8����|��V��U���u�
�
�
��}�W���&����l9��h1��*���
�
�
�
���(���&���F�C��U���u�u�u�u�w�}�W���Y���F�N��U���
�
�
�
���(�ԜY���K�X/�� ���!�4�<��'�}�(���&����l9��KN��U���u�u�u�u�w�!�(���&����l9��h1��U���u�x�u�u�w�}�W���Y���9��h1��*���u�u�u�u���(���Y���F�h1��*���_�u�u�u�z�}��������F��h��U���u�)�
�
���W���Y����l9��h1��	���u�u�u�
���(�ԶY���	��C��&���u�h�:�4�6�3��������z��Y�����d�1�"�!�w�t�W���Y���F�N��U��:�,�6�:�9��������\5��T-�����u��8�9�$�8�4�������F�N������;�u�h�8�3�����Σ�]��d��R���=�d�1�"�#�}�^���Y���F�N��U���s�:�,�6�8�3�!���Ӈ��	��Y�� ���h�}�|�n�w�}�Wϱ�����z��ON�U���;�� �!�]�}�W���6����G5��TN�U���!� ��;������*����[��_�����:�e�_�u�w�}�W���Y���F�F�����:�;��9�3�<�ϱ� ����F��
N�����9�6��6�8�}�W���s���V��^�Uʰ�1�%�:�0�$�W�W�������_��C��U���i�u��9��<�����ƣ�]��d��]���%�!�,�6�?�:�^�ԜY����R/��V��2���u�u�i�u��)�>�������]��s��<���;�}��%�#�$�ȶ�����F�-�����1�!�u�=�w�(����Ӄ��^��DN��U���!����>�)�W���������Y��U���_�u�x�4�'�-����Ӑ��@�������6�:�;�u�8�>����Ӓ��@F��o@ךU����!�u�=�#�2�����ɝ�^��U�����0�u�=�;�#�8��������`��t�����4�0�&�'�]�}�ZϪ�ӫ����R�����!�u�;�0�2�8�ϱ�Ӊ��Q	��S�Uʺ�4�4�;�0�>�1�W���DӉ��G��~F�����'�>�4�%�2���������F��V�����0�|�n�u�8�<��������bF�S��1�����&�4�;�/����	����V��T��D���:�4�4�;�9�8�^��s���%��V�����%�:�0�&�9�}����s���E��\1��3���!�;�0�%�%�>����s���E��\1�����0�u���0�����Y����[	��h�����0�9�u�#�%�1�}���T����X9��D=�����9�u��4�#�<���������X��U���!���9�3�2��������W!��Rd��Xǣ�:�>�4�&�6�<�����ƣ�R��Y=�����_�u�x�=�8��W�������Z��������'�4��w�p��������m�G����u��4�!�9�8��������X��R �����:�>��4�#�3��������\��<��\���u�2�;�'�4�0����Y�����Z������6�0�u�w�c����	����V��T��U���u�x�<�u�>�)����C����F�N�����9�6��6�8�}�W��Y����A��T�����y�u�u�x�w�3�W�������	[�=N��U����8�'�6�$�4���������Z>�����<�2�;�!�~�}�ZϷ�Yӈ��F��T��D�ߊu�u�:�!�:�-�_���Y����a��CN��U���u�u�u�u�w�}�J���5����R4��R�U���u�u�u�u�w�p��������RǻN��U���%�0�9�u�w�}�W���Y���[�x��6���u�u�u�u�w�}�W���Y�������*���<�_�u�u�w��������F�N��U���u�k�:�!�%��������F�N��U���u�;�u�:�;�<�}���Y�ƿ�[��N��U���u�u�u�u�w�}�Iϱ�����F�N��U���u�u�u�u�z�}��������GN��V�����'�,�u�u�w�.��������WF�N��U���u�h�u��#��!�������F�N��U���x�<�u�7�8�8����Y����w��e��4���0�&�3�&�#�3�J���=����V��S
�����3�0��y�w�p����,����]��v�����>�4�_�u�w�}�3���0����V/�N��U���u�u�k�:�6�<��������F�N��U���x�u�;�u�>�3���Y����G	�d��U���&�4�4�;�>�8�W���Y���F�
P��1�����'�4��}�W���Y���K�^ �����0�}�b�1� �)�W���Y�����T�� ���9�1�u�u�w�}�W��Y����F��C8�����u�u�u�u�w�}�Zϱ�ӄ��_��=N��U����6�8� ��}�W���Y���F�	N������!�y�u�w�}�W���Y���K��B����� �
�}��:�1����s���F��T��:���u�u�u�u�w�}�W���GӉ��P��B��N���u�u�u�u�w�}�Z����ƈ�G��C1�����%�0��'�]�}�Zϒ�����[��B�����'�8�!�0��8�4�������]F����ʡ�0�u�'�u�2�8��������P��=N��Xʼ�u�=�u�4�'�8��������l�G�����4�#�%�4�2�8�[�������9F��R	�����u�3�4�#�'�<����PӒ��]l�N����� ��!�4�>�����DӀ��@��N��Uʺ�6� ��!�>�8�W��Q����A�	N�����&�h�u�e�~�f�W���YӉ��P��B�����i�u�:�=�%�}�I�������[�^��\�ߊu�u�9�<�w�4��������|��t��U���;�u�u�u�z�}����Ӊ��P��B�����<�0�<�u��>����/������R��U���=�<�u�=�]�}�W���TӒ��V��[��U���9�u�<�1� �)��������@F��RN������>�!�8�9�W�W���Y����|��B������!� ��9�z����PӒ��]l�N��Uʺ�6� ��!�6�4�'���Y����r��Z!��#���1�_�u�u�w�1����Y���	��T�� ���9�1�<�0�k�}�6�������R
��g��U���:�6� ��#�<���Y����������u�u�x��#�5��������\��B�����!�8�u��4�0��������@��CךU���u�3�:�6�"���������[��N��U���:�6� ��#�4����DӉ��P��B�����u�u�u��4�0����	���F��T��:���n�u�u�u�2�9���Y����]��QUךU���u�'�6�&�l�W�W��-���� ����U���4�9�1�1�%�3�W���Y����AF��RN�����<�;�:�u��.��ԜY����]F��D�����:�u��&�#�0�Ͻ�����V��C�����u�;�!�<�w�2����Y���@��RN�����:�%�;�;�$�>����Y����V��F��%���y��:�>�6�s����P���K��RN��U���u�4�!�!�>�}��������Z��C�����<�&�"�,�#�}����/Ӡ��rl�C�����4�{�u�:�w�8��������[��^ ��U���u�;�!�<�w�2����������V��U���u� �0�!�6�}����Ӓ����V�����!�u�4�u�2�)���Y����W��U�����x�u� �4�>�3����Ӈ��@��^��Ǵ�&�'�0�u�$�>��������Q��_��#ʱ�4�'�8�_�w�p�>�������G	��RN��U���&�u�&�9�9�}�Ϫ�ӵ��C
��[�����<�0�1�9�.�}�Z�������[F��^�����0�_�u�x��)�Mϗ�Y����F��C8�����9�<�u�<�6�1�����Ƹ���R�����u�=�9�u�#�}�Z���Y���Z��E��U���;�<�u�<�;�.��������]�������&�!�1�4�$�/��ԜY���F�:��U�����u�<�0�<�W�������R��C��U���0��9�1�3�/��������F�N��U���;�u�0�%�>�}����Ӏ����[��ʺ�0�6�6�0�6�)�Ϫ�Ӡ��Z��Y�����u�&�;�7�2�(����?���]	��D;�����0�n�_�u�z�5����Y����C"��!��#���1�9�%�u�z�+����Ӎ��@��V��E�ߊu�x�=�:��}�%���Ӈ��u��e�����x�#�:�>�6�>�ϭ�����|��B�����x�=�:�
�w�1�W���	����Xl�C�����4�6�u�:�$�9����Q����F��C8�����%�|�u�x�!�2�����ƿ�P��x������9�u��#�<��������]��NN������:��%��)�^���YӁ��V����U�ߊu�u�u��$�)����G����F�N��Uʦ�1�9�2�6�m�}�G�ԜY�Ƽ�A��V�����u�u��&�#�`�W���?����V��N��U���u�u�u�u�w�}�W��Y���Q	��R��U���u�6�;�u�w�c��������G��q(�U���u�u�u�u�w�}�W������\	��V ךU���u�9�u�u�j�}��������F�N��U���u�u�u�u�w�}�Z����ƿ�W9��P��U���u�6�u�u�w�c��������Z��v������9�1�<�2�q�W������G��X	�����u�u��u�w�`�W�������G0��^
����u�u�u�u�w�}�W��Y����@��[����u��&�!�6�W�Wϙ�����V"��V!��O���3�'��6�9�8�W�������_��R�����d�1�"�!�w�}������ƹF��R ����� �%�!�4�6��M���YӀ����YN�����6�8� ��1�_���0����A��P�����4�0�u�u�w�p��������u
��s��:��� ��!��8��W���Y����[	��h��'���!�4�u�e�]�}�W���T����X9��V<�������2��$�)�W���Y����[	��h��0����4�9��#�(�1�ԜY���K��X��ʖ�>��8�9��6�W���Y����[	��h��1ʺ�6� ��!�>�8�_���0����N��=N��U���x�=�:�
�w�����������=��<���-�}�|�u�w�}�8�������R ��G'����!�u�:�>��1����Y۔��l�N��Uʲ�;�'�6�8�'�u�W���Y�����D�����k�r�r�u�z�}��������T��S��E�ߊu�u�u�u�8�)����Q���F�N��'���!�h�u���:�%������F�N��U���u�x�u�;�w�2����s���F�N�����u�k�&�;�5�8�������F�N��U���u�x�<�u�5�2����Y���F�-��U���h�u�4�%�2�1�[���Y���F�N��U���x�u�;�u�#�����s���F�N��U���u�k�:�6�"������Ο�P/��R�����u�x�<�u�$�9�������F�N��$���u�h�u��4�0�����Ο�P/��R�����u�x�u� �w�)�(���������D���ߠu�u�u�x�!�2����=����w��x�� ���!��:��w�}�W������l��e�����u�e�_�u�w�}�Z�������R4��R��9���2��&�!�w�}�W������l��r ��0���9��!� ��W�W���Y�˺�\	��VN��ʆ�8�9��>�w�}�W������l��sN������!�<�0��-�>����Υ�9F�N��X���:�
�u��$�>��������5��~ �����|�u�u�u��)��������C7��R �����:�>��9�'�.�WǬ����F�N�����6�8�%�}�w�}�W���YӍ��@��V��K��r�u�x�u�9�}��������	[�IךU���u�u�:�!�:�-�_���Y���F��e����u���2��.����Y���F�N��U���u�;�u�:�;�<�}���Y���F��YN��U��&�;�7�0�"�-����Y���F�N��U���<�u�7�:�2�3�W���Y���%��N��H���4�%�0�9�{�}�W���Y���F�N��X���;�u�!�
�8�4�}���Y���F��N��U��:�6� ��#�4����	����V�^G�U���<�u�&�1�;�:����Y���F��fN��U��u��6�8�"�����	����V�^G�U���u� �u�!��2����DӍ��@��VךU���;�u�0�0�6�8�0�������F��C*�����n�u�0�1�0�3����Y����A��s��:���_�u�x�u�$�4�Ϫ�Ӏ��R
��X����� �&�u�&�4�(�8�������[��X1�����;�&�6� ��)����5���9F��v������i�u��4�0������ƹ��T�� ���i�u��6�:�(�;���B���WF��{U�