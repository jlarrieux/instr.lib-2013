-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����X��b�����&�#�1�x�w�(����Y����$��[�����u� �&�4�#�<�W�������A	��t��ʖ�;�4�_�x��4����Y����V��-��;����&�<�2�z�}����Y�ƃ�G	��EN�E�߇x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T����F��]�����<�=�u�4�>�3�ϗ�
����V��-�����!�:�_�x��1�%����ƞ�@��R
חXʛ�!�:�4�u�9�)�����ƅ�G��V�����8�!�:�_�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���x�x�u� �'�.�M���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W��T�Ɯ�T(��C�����u�<�9�%�8�4�ϭ��Ư�^��[�����1�3�;�!�8�.����Y����]	��N����%�:�<�0�w�$�>���Y����R��N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�z�W�Z���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���K��C�����,�0��:�2�3����ӏ��@	��V��U���8�!�=�!�2��W����ƫ�Z��^ ��U���u�u�x�x�w�(��������\��X�������&�0�w�4����������V
�����u�u�,�0�5�)�W���Y��ƴF��RN�����&�9�>�9�w�2�����Ƹ�VF��^�������%�!�2�3�W�������E��X�U���_�x��'�9�0�W���^�Ư�_
��RN�����=�!�3�!�%�}����
����\	��V �����w�<�u�u�w�}�Z�ԑTӖ��Q��NN�����u�=�<�0�1�/����Y����\��[��U���u�u�u�u�w�}�W���Y���F�C�X���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�z�p�W���Y����V��X �����0�;�7�:�2�3����
����\����U���!�:�0�&�6�}����Y���KǶN��Rʼ�u�:�u�;�!�/����Y����A��X
��ʸ�4�u�!� �u�}�$���Ӈ��Z��_��U���u�x�_�x�;�:�Ϸ�Y������Z�����u�6�<�0�;�*�W�������V��XN�����=�u�u�u�w�}�W���T�����^�����u�:�#�'�>�3�W���Y������G��U���0�u�!�
�8�1�������F�N��U���x�u�!�
�#�����W�Ƙ�VF��C��X���u�0�&�:�$�(�Ϫ�ӑ��W��V��U���u�u�u�u�w�}�Z��Yђ��q	��R�����0�:�w�u��(����Ӗ��U��C�����!�!�0�!�2�<����T����F�CחXʧ�&�9�&�7�#���������@����U���<�0�9�"�4�3�����ƿ�]��C�����;�u�u�x�]�p��������K��T��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���l�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�x�x�u�9�)�Ϯ�
������@�����w�0�<�0�w�(�����ƪ�AF��S1�����#�6�:�u�?�)�W���T���R��[��U���u� �0�<��)�W�������F��^����� �&�2�0�y�}����
����V��N��X�߇x�<�u�0�<�.����
����\��h�����<�u�:�u�;�<�Ͽ�Y����T�������;�8�0�{�w�p�}��.�ƣ�G��@��U���/�'�u�4�w�3����������C��U���9�3�y�:�w�<�������F�d�U���!�0�8�1�;�s�W���Y����U��C�����0�:�w�4�3�����Y����Z��Y
��U���u�u�u�x�z�}����Y������U��Yʰ�%�6�4�9�w�5�Ͻ�����TF��V
�����0�<�!�'�w�4����Y���9K�D��U���&�1�7�!�m�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���x�_�x�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W��s����Z��[N������!�u�u�#�����&����\�N�����u�|�u�u�w�}�W���Y���F�N��X���u�{�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�p�Z�������w��R��/���&�d�|�s��)��������F�*��'���0�!�s��2�;��������F�=C�U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�x�_�z�����
ӏ��V��SN��U���%�"�<�0�%�p����Ӆ��C	��Y��U���6�u� �u�?�}�W���Y���K��O�����:�8�;�u�!�/����5����U��C��U���!�0�%�6�6�8����W���F�N��U���x�x�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W��T�ƅ�G��\N��ʆ�4�9�'�4�3�����Y����G��DN�����'�4�:�4�;�}�Ͻ�����~��N����4�1��-�w���������_�C�����!�:�u�4�2��Ͻ�����@F��C�����8�;�u�u�z�W�Z�������@O��R�����;����6�9��������VH�c�����u�<�u� �4�4�������K��C�� ���7�u�4�9�3�����������^ ��:����2�<�!�;�)��������O�N��U���u�u�x�x�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y���F�N��U���u�u�u�u�w�}�W���Y��ƴK�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���_�<�'�'�w��2�ԜY����z#����*���<�
�d�a�6�1�}���
�ƅ�v#��B�����!�{�9�n�]�<����Y����Z3��[�����&�_�u�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��s���3��Q�����,�!�%�&�w�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���9l�C��U���9�4��6�8�}�Ͽ������B��U���2�i�u�u�1�?�������G��'������6�:�u�$�<����Qӈ��F�������k�u�3�<�#�:��ԜY����(��B��#���:�u�&�4�%�$�_ϰ�������P��K���3�;�!�'�;�W�W���ӵ�� T��N1�����'�4�u�u�6�(��������X������9�2�6�#�4�2�_������\F��d�����u�9�d��.�)��������F��C��ʧ�;�0�i�u�w�;��������l��C��D���:�;�:�e�l�W�W��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K��N�U���0��;�0�$�2�W�������@l�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�_�u�z�<����Y������A�����u�d�u�k�#�(�}�������\��X1�����;�}�u�u�#������ƾ�G�������n�_�u�x�6�)�����Ư�]��D��Y��r�x�u�'�2�}��������G	��X�����!�#��"��}�W���&����Z�E�����:�9�4�n�]�}�ZϿ�����[�������<�;�u�d�u�p�WǪ�����R
��d�����!�:�u�:��2�����������*���<�
�0�!�%�}����Ӥ��_��a����_�u�x�4�#�+�W���Ӆ��E��^��U��w�x�u�3�;�8�W������U��C��U����:�0�;�2�)��������DN��N�����2�6�#�6�8�t�W���Y���F�N��U���u�u�u�u�w�}�W�������]F��X�����!�'�_�u�z�}����ӎ��[F��Y�����y�!� �u�i�z�P�������Z	��C�����2�6�7�o�5�2����Y����A��C
�����6�_�u�x�w�>��������\��E�����4�&�u�k�p�z�Wϸ�����]F��h=��9���6�6�<�0�8�u�W�������]O��R��ʦ�1� �:�<�l�W�W������VF��P�����'�<�;�u�#�(�[ϸ����X�^��Uʳ�;�!�:�u�8���������G	��UN�7���0�;�0�!�%�}����ӕ��l
��^�����'�_�u�x�w�>��������P	��R�����}�'�0�u�6�.�^��Y����9F��B �����!�
�!��0�>��������E��@F��Oʗ�:�0�;�0�#�/�}���Y���F�N��U���u�u�u�u�w�}�W���YӔ��F��D�����6�#�6�:�l�W�W��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K��N�U���6�3�;�!�8�.�W��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�=d��X���0� �;�u�w�)�(�������P����ʙ�;�!�u�<�$�}�����Ƹ�A��=N�� ���<�;��'�$�����Y�Ƣ�G��[G�����;�&�1�9�0�>������ƓF��� ���u�u�!�
�8�4�(�������Z��{�����<�&�u�9�w�8�W���^��ƹ ��T��ʚ�0�}�0�2�?�g�������A��E �����:�<�
�0�#�/�}���T�ƾ�G��DN�����2�:�u�4�2�o��������9F��B ������2�}�'�w�}�������A��E �����4�n�_�u�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K��^��6���4�<�:�u�"�>����s���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X�ߊu�x�'�!�%�.��������AF����U���u�;� �&�w�;�����ƀ�A����U���;�0�0�|�%�)��������A]ǑN�U���u�&�?�&�w�3����Y����G	��V��9���0�{�u�x�w�1����
ӈ����G�����,��;�9�4�)�W���s���3��X�����=�u�9�4�w�8��������Z��_�� ���0�u�x�4�>�.�:����ƀ�A��5�����'�u�;�0�2�}����ӏ��V��jUװU���u�0� �;�w�5�W�������\ ��_�����;� �&�u�1�3����Y����_��VB��Oʼ�!�2�'�u�2�(�Ϸ�����lǻC�8���<�u�;�!�2�}����Ӆ��_F��V������"�#�'�w�5�Ͻ�����+��N�� ���x�u� �!�"�8��������W��Y��UȂ��{�>���4����
ݫ����L��ʴ�:�1�u�x�w�2��������Z��C�����0�<�!�:�w�2�Wͳ�����F��Q��ʼ�_�u�x����������p��^ ��&���9�'�<�u�%�?����
����V�N�U���4�u�&�;�#�.��������JF��Y�����u�{�_�u�z���������[��[��U���9�'�!�:�w�3��������Vl�C������;�<�u�:�1��������V�^ �����'�!�'�u�9�8����s���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X�ߊu�x��6�8�}����Ӏ��P��YךU���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�]�}�Z�������U��C��ʧ�!�'�u�=�w��Uϱ�Y����JF��CN��U���u�0�!�'�'�.��������F��^��:���6�:�u�4�0�g��������l��C��U��� �;�&�1�"�2���YӀ��P��YN��#���:�u�4�2�m�(��������V��YN�����:�<�n�u�1�3����Y����P��F�����:�0�;�2�)����������[��N�ߊu�x��0�2�;��������V��YN������w�:�u�!�/�W���Y����[��R��ʥ�&�0�u�;�w�;�����ƍ�W0��C��]���u�u�!�
�8�4�(������A��E �����9�2�6�_�w�(����ӧ��e��X�����o� �&�2�2�t�����ƿ�W9��X	��N���3�;�!�:�w�3�!�������A�,������6�:�|�%�)��������]]ǑN�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�u�z�}��������J��R��U���'�7�!�&�w�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���9l�V�����0�&�;�=�2�}�W�������F��C�� ���&�;�7�4�<�?�������R��N����� �0�&�;�2�>����Y�ƿ�A��d�����<� �0�&�9�8��������]������_�u�!�'�5�)�W���&����\��X����u�4�!�<�"�8��������G9��V��U���:�9�4�n�w�<��������J��V����<�!�2�'�]�}��������K��E��U���!�<�2�_�w�)�����ƿ�]9��T�����u�u�:�9�6�f�WϿ�����G��X�����u�u�!�<�0�W�W�������VF��Y1�����7�0�u�u�8�1���s���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�u��;�#�2�ϸ�ӕ��G����ų�0�1�u�<�?�3�Ϩ�����F�N��ʺ�u�=�&�u�"�>����Y����A����*���<�
�0�!�%�*����Y����VF��=N��X���x�u�:�;�8�m�[ϩ�������V��ʡ�u�g�<�u�#�4�W���Y����Z ��S@ךU���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�]�}�Z�������V��N����x��!�'�w�}�E¼�Ӑ��G	��@��U���&�`�u�c�w�3�W��
��ƹK�\8��F���h��!�<�$�u�[��U����]ǻC�U���u�:�<�0�#�<�W���Y����A��V��ʸ�&�u�0�0�4�2����Ӗ��V��R��Yʦ�u�:�_�u�z�0��������\��RN�����u�=�;�,�"�>��������@H���R���;�!�0�u�6�}����T�ƫ�GF��RN�����0� �!�!�6�}����Y�����������3�'�!�0�2�)�Ϯ�����F���ʶ�0�'�_�u�z�6���Y����V��C�����0�h�}�y�f�q�F���B���l�C�����;�4�c�x�>�}����ӑ��[F��C��Y��u�y�4�1�a�}��ԜY����e��N�U����!�}�g�w�q�A���J���O��N�U���9�0�;�!�!�1�}���TӍ��PP��S�����!�}�;�<�2�`�_��M����P��N��K��n�u�x�_�w�p�%����ƭ� T��^�����'�"�!�u�>�}�W���s�����T]�I���0��!�f�l�}�Z�ԜY����V��YN��F���<�u�0�!�%�*�����Ƨ�\��CN�����u�;�!�0�!�1�ϱ�Y�ƿ�T�������-�:�_�u�z�<�ϼ�Ӎ��V$�������:�u�=�u�6�(�W���ӕ��]��T������0�u�x�w����E�Ɵ�G$�������y�-�:�|�8�}����ۍ��V$��N�����_�u�x�u�z�}����Ӈ�K��CN�����u�=�'�u�>�}�5����ƿ�GF����ʴ�1�!�0�-�8���������AF��=N��Xʴ�&�2�0�u�8�)�ϼ��ƿ�R��Y	��ʷ�!�>�:�_�w�p����J���5��u������!�u��5�}�ύ�����WN��X�����0�1�n�w�p�}���TӨ��VF��V��?���<�9�u�4�w�8��������AJ��YN�����0�y�:�u�w�)�(�������P��d��X�ߊu�x��!�$�.�ϩ�Y������R�����'�2�&�0�y�}����
Ӓ��	����U���1�u�!�_�w�p�W��Y����V��������0�<�9�{�0�������F����ߊu�x�u�8�2�n�W��Q����A�	N��R��u�x�u�u�1���������+��R	����:�!�;�u�?�3�W��Y���^0��\��7���<�|�i�u��?�}���T�����T]�����0�1�&�w�2��������Z��N�U���0�<�9�n�w�p�W����ƥ�l�C�����'�6�&�n�w�p�}���Tӧ����RI�����;�"�"�,�]�}�Z���T�ơ�V��R��&���<�}��7�>�q����PӉ��`��^��]���0�<�9�y�:�2�1������K�N��U���u�u�"�0�w�8�$�������~��PB��<���'��|�0�$�}�������A��UךU���u�x�u�=�$�}��������R��V��U���3�9�<�u�2�)�����ƻ�V��E�����;�u�0�1�9�W�W������G��N�����1�'�!�0�8�9� ���s���9F�N�����h�}�!�0�$�`�W��P���K��V�����|�o�u�d�l�}�Z�������y	��^��8���1�"�!�u��8����P���F�N��U���u�u�h�&�3�1��������AN��h;�����1�d�y��2�4�������9F�N�����:�:�!���:�W�����ƹK��N�U���u�:�u�=�w�8�W���C���l�C�������'�}�.�8�[ύ�����X$��N��U����0�1�>�8�����Y���lǻ�����;��!�<�$�����
����R��V�����n��o�;�#�/���Y���A��E �����:�<�
�0�#�/�}�������\��R���1�-�o�;�#�/��ԜY���F�N��U����9�o�&�3�1����C���]ǻN��U���u�u�u�u�w�}�W�������	[�G�����;�&�1�9�0�>������ƹ ��T��ʆ�!�<�}�;�2�}�W�������1� �� ���u�h�f�|�%�)��������T��A����u�3�;�!�8�}����ۯ��V� �� ���n�u�u�u�w�}�W���Y����R
������n�u�u�u�w�}�W���Y����\��V�����h�f�|�'�#�/�W���&����P9��T��N���3�;�!�:�w�8�1���ۯ��V� �� ���n�u�u�u�w�}�W���Y���0��T�����;�1�_�u�w�}�W���Y���F�`N����'�9�o�u�e�}����ӕ��l
��^�����'�_�u� �4�4�ύ�����WN��S��Oʻ�!�'�9�_�w�}�W���Y���F�N����&�1�9�2�4�+����B���F�N��U���u�u�u�u�w�<����Y���O��R��ʦ�1�9�2�6�!�>���YӀ��P��YN�����9�}�;�0�w�}������ƹF�N��U���u�u�u�u�6�}�W�������9F�N��U���u�u�u�u�w�}�W�������	[�G�����;�&�1�9�0�>������ƓV��g������2�<�!�;�)���s����R��U��U���� �<�<�>�.��ԶY���g��Z��U���4�0�,�:�w�5�W�������AF��G�����!�:�&�<�w�2� ���Ӊ��9F�N��U���u� �6�<�9�}��������VF��RN�����:�{�u�9�w�5�W����ƪ�]��X ��U���u�0�<�0�#�8�ϼ�����AF�������u�=�u�4�2�;�������F�=N��Xʜ�u�=�&�6�$�q��������]F��SN��*����2�6�4�2�)�ϼ�
�ƪ�]��X �����x��0�#�4�2�W�������A��^��ʶ�9�u�=�u�6�8����������E�����{�u�x�u�?�}����ފ����A�����8�'�9�u�9�8�Ϫ�Ӕ��F
�������7�&�_�u�z�;�������F�=N��Xʁ�<�u�%�'�6�5��������A��T�����4�:�;�u�1�>�������GF��DךU���6�;�0�!�6�8�W���Y����E����ʴ�&�4�9�%�6�8�Wϗ�Y����@��[���ߊu�x�6�;�2�)�����Ư�A��CB�����7�2�u�;�#�8�����Ư�]��C��U���_�u�x�4�:�.�W�������V��XN�����u�:�!�0�>�8����ӄ���������x�6�;�0�$�2�Ϫ�����E��=d��X���0�<�0�!�2�?��������@��=N��Xʀ�9�>�u�=�w��2Ϻ�����	l�C��U���6�<�;�!��4�_���Y����_	��TU�����o�7�!�u�2�(�ϼ����K��B�����'�0�u�:�$�3�Ͽ�����]��X �����!�:�u�:�w�5�W���ӑ��]l�C�����;� �u�4�w�}��������F��X�� ���y�"�r�0�0�8����Y����V��N@ךU���6�<�;�!��2����Yە���h�����u�0� �;�5�2�������Q��Yd��Uʧ�!�'�u���m�_���^���9F��Y
�����:�0�;�_�w�p�W�������\��E��U���0�u�;�4�w�%����Ӊ��A��EN�����|�u�3�;�#�2�W���;����R��C��9���}�u�u�!��1����Y����A��X�����&�u�7�2�9�}�WϬ�����2��o^���e�|�_�u�9�}��������r��A���ߠu�x�u�u�2�4����Ӆ��E��R�����u�=�u�4�2�>������ƹ ��T��ʡ�
�:�9�4��>����Y�ƿ�W9��P�����:�|�'�!�%�}��������G	��^ךU���4�<�7�0�%�<�W�������]0��C��ͧ�;�0�n�u�5�:����YӀ����YN�����4�2�u�:�'�}�W�������ZO�
N��*���9�4�}�}�~�f�W�������\	��=N��U��� �;�'�4�l�}��������\
��Y8�����_�u�x�u�w�8��������\��E��U���;�u�;�0�>�)����	����\� ��W�ߊu� �6�<�9�)�(�������V��E/�����:�}�u�u�#�����&����\�N��U���u�u�u�u�w�}�W���Y���F�N�����'�u�:�9�6�����Y��ƹF��V�����'�4�u�u�8�1��������@A��Y	��N���7�2�;�u�w�;�Ϸ��ƾ�R
��V ��U���%�u�u�u�%�<�_���C�Ƹ�l$��[��4���#��"�&�>�t�}���Y����_	��d��Uʧ�!�'�u�#�;�W�W���Y����\	��V ������!�#�� �W�W��Y����Q�������<�;�u�3�9�)��������	��TF��Oʷ�:�0�;�u�2�(�ϭ�����T��^ךU���<�_�u�u�1�?����s���F��C��U��n�u�u�0�$�W�W���Y����A�I�U���0�1�<�n�w�8�Ϫ�&����\��dךU���6�<�;�!��)�;�������E��@F��Oʷ�:�0�;�u�2�(�ϭ�����T��^ךU���<�_�u�u�2�(�ϰ�Ӓ��`��X	��]���_�u�;�u�8���������Z��X���� �6�<�;�#���������P����U���9�4��6�8�t�����ƿ�W9��P�����:�u�&�u�w�+�����ƾ�R
���*���<�
�0�!�%�?������ƹ��^ ךU���:�u�u�;�%�<�P����Ơ�\ǻN��U���9�<�u�h�#����������d��Uʰ�1�9�:�n�w�}�����ƾ�R
��N��ʡ�
�!��2�4�8����s����F��^�����!��2�6�2�)��������DN��N�����;�0�!�'�]�}�W���Y���F�N��U���u�u�u�u�w�}�WϬ�����@��[�����6�:�u�&�w�?����Y����V��YN��ʡ�
�!��2�4�8������ƹ����&���:�<��6�8�����5����9F��B ������'�&��9�)�W�������_O��R��ʦ�1�9�2�6�!�>����
�����^��ʃ�6�u�!�
�8�4�(��������{�����o�u�:�=�%�}�I���^��ƹ��^ ךU���0� �;��4�W�W���Y����@]ǑN�����:�u�;�&��3����Y����A���� ���&�1�9�2�4�+����Y��ƹF��V������6�u�!��2��������W��XN�����|�o�u�:�?�/�W���^���9F��R	�����u�0� �;��>�}����ƃ�V��=N��Xʙ�2�u�0� �9�}��������TF�������g�9�2�'�#�0�Wϛ�������[�����o�u�x�_�w�p�����ơ�KF��=N��X���2�;�'�6�]�}�Z���Yӑ��G������u�h�f�_�w�p�W���s���F��X�����x�u�u��9�g��������T��A�����<�!�x�u�8�3���B���F�N����<�u�;�<�9�9����Q����[O�
�����e�n�u�x�w�}�W�������F��C
�����_�u�x�u�~�W�W������F��N�����:�u�:�g��:�MϮ�
����VO��R��ʻ�!�'�9�<�]�}�W�������4��B�����u�4� �4�l�}�WϨ�����VF��^�����u�u�4� �6�f�Wϼ���ƹF��R�����u�h�e�_�w�}��������\�v��D�ߠu�u�"�<�2���������F��[�����u�u�=�3�2����Y����G��E	��U��u�u�u��#�/�!���C�ƞ�G��a��^��_�u�u�;�w�2��ԶY����V��YN������9�_�u�9�}���s����F��^��9���0�}�y�u�w�3����PӔ��F��^ �����<�_�u�0�>�W�W���Ӈ���_��U���u�'�!�'�w�f�W�������F�N�����u�n�u�u�2�9���YӃ��*��P�����3�;�!�:�w�0����Q�ʮ�	F��C�����0� �;�<�#�:�Ϸ�s�Ʈ�T��N�����u�u�u�=�9�}�W�������]F��=N��U���0�u�u�u�%�)����B����������;�u�8�9�2�f�}���TӲ��@��B �����u�0� �;�#�8�U���Y����E����U���!�0�#�6�8�}����ӏ��F��Y�����'�0�!�'��/�W�������T��A�����'�!�'�u�#�����ӏ��F�A�����u�0� �;�6�}�W���&����Z��N�����u�u��!�%����Y���9F���U���;�4�2�'�9�8����s���F��C��#���o�u�0� �9�<�W�������]ǻN�����:�%�_�u�w�8����+����]0��d�������6�:�l�W�W�������)��R�����'�u�u�;�>�3����������h�����<�_�u�0�>�W�W�������)��R��¦�1�9�2�6�!�>�������9F��Y
�����!�'�_�u�1�3����Y����P��F�����:�0�;�2�)����������[��U���u�7�2�;�w�}�����Ƙ�l$��[��]���0�!�'���)�;�������\��E	��\�ߊu�;�u�'�2�)��ԶY���g��RN�����:�&�'�!�%�}����8���\ ��A��U���u�3�!�0�!�>����������N�����:�u�;��4�2�Wǿ�����G��X	��*���!�'�u�0�"�3��������PF��=N��U���<�7�0��#�/�!���Cӕ��l��P�����0�<�_�u�w�8��������A��d��Uʳ�'�<�<�u�%�z����Y����9F�N�����;�4�u�h��)����Ӈ��������u�;�u�:�'�W�W�������4��B����u�0�1��3�8����s����F��^��4���0�!�'�}�%�}�W�������F��C��U���
�9�2�6�>�W�W������F��C��U����6�:�}�#�����&����\��E	��N���0�1��1�2�)��ԶYӀ��P��YN�����!�'�}�'�w�}��������G	���� ���7�:�0�;�>�W�W������F��C��U����:�0�;��9����۲��`��X	��#���:�}�'�|�~�W�W���Y����V��EUװ���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�W��?����Z	����U���!�;�u�<�$�<�ϼ�����W��^��ʴ�#�6�:�_�w�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���9F�N�����&�4�&�1�;�:��������D����U���&�6�'�0�'�3�����ƅ�W��DN���ߊu� �6�<�9�����
ۯ��Z��T�����4��6�:�l�
�Mϰ�����\�\�����'�u�!�
�8�4�(�������@l�N�����9�u�4�4�m�.��������V��EF��Dʱ�"�!�u�|�]�}����s���w��T��]���0�&�h�u�g�t�}���Y����ZF��'�����r�4�2�u�8�-�W���YӢ��RN��S��¼�|�o�u�d�l�}�Wϻ�ӊ��C]ǻN�����;��!�n�w�8�ϸ�����]F��C,���ߠu�x�u�0�"�3�W�������T��A�����<�=�7�!��9�����Ƹ�5��=N�� ���<�;��!�>�u����Y�Ƣ�G��[UךU���u�u�u�u�w�}�W���Y�ƿ�W9��P��O���d�n�u�u�w�}�W���Y���1� �� ���u�h�f�|�%�)��������T��A�����&�u�u�#�%�<���������h�����0�!�'��f�9� ���Y����F��P��U���x�&�;�=�$�.����
����l	��=N��U���0�!��1�/�a� Ϭ�	����/��R�� ���7�u�0�&�#�<�W���
����Z��R���ߊu�u�x�,�#�8��������R��X ךU���4�4�o�u�8�5����G����]ǻN������1�-�u�j���ԜY�ƾ�G��*���ߊu�;�u� �4�4�ύ�����9l�C�����;�u�u�!��2����������_N��ʷ�!�6�'�0�'�3�����ƅ�W��D����� �6�<�;��)��������	F��C�����u�u�4� �6�}�J��PӔ��F��D�����6�#�6�:�w�.�Wϼ���ƹF��R��ʆ�!�<�}�;�2�`�>����ƚ�_[�I�"���|�_�u�;�w�(����ӵ��q��=d��X���0� �;�u�w�)�(�������P����ʷ�!��1�-�w�8�W���*��ƹ ��T��ʆ�!�<�}�;�2�}�W�������9F�N��U���u�u�u�u�6�}�W�������9F�N��U���u�u�u�u�w�}��������U���� ���&�1�9�2�4�+����Y��ƹ��^ ךU���0� �;��#�4�_�������]��N�����:��1�:�>�u����Y����]ǻ��U���6�<�;��#�4�L�ԜY����V��Y��U���
�:�<�
�2�)�Ϫ��Ƥ�@F��[N�����0�u�!�u�z�}�����Ƽ�@��X �����4�0�u�,��9��ԜY����G��=��3���1��1�-�m�3�������F�N��U���u�u�u��;�g��������9F�N��U���u�u�u�u�w�}�W�������	[�G�����;�&�1�9�0�>�����ƥ�9F������0��!�u�w�)�(�������P��9��U���;�:�e�u�j�u����
���V�d�����;�u�u�x�$�3����
Ӓ��]��C���ߊu�u�&�0�#�����Eӱ��V��CN�����u� �!�7�w�8�Ϫ��ƛ���R��ʰ�'�'�_�u�w�.����Q����_��C��U���0�|�i�u�]�}�W�������D��[N��U���u�<�u�:�1�)��������F��A�����'�:�n�u�w�p����������Y�����;�u�u��#�u�Z�������/��R��O���!�
�:�<��8��������VN��[B��X���0�|�n�u�w�/����Y����l�R �����!�:�u�0��8��ԶY���a��E ��ʦ�1�9�2�6�!�>��������R��V�����;�1�4�_�w�p��������\��^�����6�!�1�7�w�3���YӀ��P��YN�����9�}�;�0�w�}������ƹF�N��U���u�u�u�u�6�}�W���&����P9��T��N���u�u�u�u�w�}�W���Yӱ���B��U��f�|�'�!�%�}��������E��X�����7�2�;�u�w�/����Y����Z��'�����1�-�u�6�`��������e��N��K���_�u�;�u�"�>����*����V
��=d��X���0� �;�u�w�)�(�������P����ʽ�&��9�'�#�/�������F��RN��ʥ�&�!�:�u�9�4����Y����]��d�����!�:�u�0��8�Ǘ������B��N���u�u�u�u�w�}�W���YӰ��\��V����u�u�u�u�w�}�W���Y����\��V�����h�f�|�'�#�/�W���&����P9��T��U���u�7�2�;�w�}�����Ɵ�G ��[
�����h��1�-�w�<�Jъ�&����T��8��Yʂ��1�-�y� �c�^�ԜY����U��C��U����0�1�_�2�9�'�������\��g�����9�!�0�n�]