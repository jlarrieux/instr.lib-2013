-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����B"��V#�����#�1�x�u�"�5�����Ǝ�X��C�����;�9��:�2�)�W�������4ǶN����g�u�0�0�5�/�E��s��ƴK�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���_�x�}�|�e�l�W��� ����GF��C�����;�!� �0�#�}��������]l�/��U���=�&��&�%�8�}��7����]��~ �����;�&��!�%�<�W�������Z	��C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�]�p�'�������g�������;�u�8�9�:�3�Ͽ�H�Ʈ�GJ��GN��U���0�%�u��z�<����T���@��CN�����0�{�u�=�w�.����<�ƿ�T����ʶ�;�'�9�u�%�)��������\F��Rd�U����y�;�!�#�8�����Ɗ�l�=C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�_�]�4����Y����l�B�����{�!�
�:�>��F������F��RN����� �0�<�
�#�s���s����J��R��U���;�9�!�
�1�W�����Ɣ�_��t��9���_�<�'�'�w��$���s����f(��~#�����:�0�!�{��f�Z��� ����@��C�����0�:�_�_�9�4�ϛ�=����V��NN��U���:�!�_�u�6�-����J���	F����*���<�n�u�&��)�>���Y�����D�����6�#�6�:��j��������l�D�����;�u�u�o�>�}��������9F��D/�����u�u�u�u�9�.��������V��EF����!�u�|�_�w�.�������F��X�����9�2�6�#�4�2�_������\F��G������!��:�/�L�Զ����G��B��'���:�u�$�4�6�8������ƹ��G�������g�_�w�}����Q���F��[��U���&�1�9�2�4�g�W��B���F��T��ʦ�1�9�2�6�m�}�G��Y�����N��U���
�:�<�u�j�z�P�ԜY���RF��^ �����:�<�
�0�#�/�CϺ�����O��N��Uʤ�o�:�!�&�3�1����s���F��N����&�1�9�2�4�f�Wϻ�Ӆ��C	��Y�U���#�:�>�&�0�)��ԜY�˺�\	��D���ߠu�&�2�4�w�.����
����_F��D�����6�#�6�:��}�������9F��^	��ʦ��!��!�8�?�Mϭ�����Z��R����u�:�;�:�g�f�Wϭ�����@��C�����u�o�&�1�;�:��������Q��X����u�h�}�!�2�.�I��P����V��=d�����1�0�&� �;�a�W��I���@��S���ߠu��;��$�W�W���Y�ƥ�V��XN�U���0�4�0�u�w�p����ӵ��pU��=N��U���=�:�
�u�;�}��������Kl�N����>�4�1�&��)�>���P���K��_��*���0�&��<�2�3�W���Tސ��\�������'�&��9�]�}�W�������RF��D�����!�:�7��]�}�W�������RF��N���ߊu�u���e�%�W���:�ԉ�F�N�����4�u�_�u�w�}�W���Y����R��R-��F���u�u�u�x�w�3�W���&����PF��I����u�u�u�u�w�c��������zO�N��U���u�;�u�!��2����D����9F�N��U���u�k�&��>�8����Y���F���U���
�:�<�u�j�z�P���Y����S����1�0�&� �;�}�W���Tӏ����h�����0�!�'�a�3�*����P���F���U��&��!��#�2�Ǘ�U���	����*���<�_�u�u�w�}�D���GӉ��]O��N��U���u�u�x�u�"�}��������F��SN�����!�u�0���f�}�������U\ǻ�����}�4�%�0�;�n�^�������9F������;�
�1�0��0�������G��=N��U���&�4�4� ��1�K���
����|��X�����u�;�u�3�]�}��������@F��Y���ߠu�&��!��)�K���
����|��T����u��n�