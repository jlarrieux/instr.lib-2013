-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����B5��P�����'�#�1�x�w�(����Y����q��Ed�U���2�;�9��8�8����!����R��=C�1���o�g�u�0�2�?���H���9K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�_�x�}�~�o�F�������T��y�����u�;�!� �2�)�W���	����Z	��C�����<�=�&��$�/��ԑTӨ��Z	��[N�����8�;�&��#�/��������R��Yd�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�Zώ�����	F��^�����;�;�u�!�>�:�W���������B��ʺ�u�$�4�f�p�}�ϳ��ƭ�K��������3�9�2�s�W���Y����P��RN��ʡ�<�u�<�!�%�4�Wͭ��˼�A��R��U���_�x�u�<�w�8�ϭ�������q�����x�u�;�!�2�����Y����V�*��U���'�2�<�1�]�p�W�������C��N�����4�;�1�3�2�8����
Ӓ��GF������6�0�3�6�2�)�W���s���"��V��]���8�!�=�!�2�n�W�������X��@חX���u�u�=�&�3�.����
���� ��V��&��u�!�!�0�2�9��������Z���� ���4�:�{�x�w�}��������J	��T��ʧ�%�4�0�!�2�;����=������_N�����0�4�6�8�;�)�������F�������<�2�!�u�6�8����ӊ��Z��CN��ʶ�&�u�3�4�w�9��������`6��N���߇x�u�!�0�6�9�ϼ�����	��^�����u�<�<�2�]�p�Z���Y����_F��G�����0�4�u�&�o�>����W���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�_�9�7�6�$����B����@��R�����9�2�6�d�a�s���Yӓ����R@�����6�&�1�4�;�W�Z��� ����@��C�����0�:�3��5�<�φ�����\��^����4�,� ���f����,����~H��X�����&���_�z�.����
����A��[��*���_�0�!�!�w�,��������V��DN�����}�u��8�;�����Y���	F����*���<�n�u��:�1�4������F��^ �����:�<�n�u�$�4����6����G ��N��U���
�:�<�n�]�}�4���5����F�N��U���&�1�9�2�4�W�W�������F�N��U���;�&�1�9�0�>�}���:����Z�N��U���u�;�&�1�;�:��������Q��X����n�_�u��#��������\��YN�����2�6�_�u��)�>���Y���F������9�2�6�#�4�2�_������\F��d�����4� �u�u�w�}�W����ƿ�W9��P�����:�}�b�1� �)�W���s�ƿ�R��V��:���u�u�u� �w�)�(������9��+�����0�<�!�'�]�W��������A��c"��ʐ��;�9��;�8�W���s���E��\1�����'�_�u�<�9�1��������F��P ��]���:�;�:�e�l�}�����ƿ�`��[����0�;�_�u�z�5��������9l�C�����6�;�!�;�w�2����
ӎ����NN��6���4�1�!� �w�2�W��� Ӓ��@J��E��ʡ�0�u�x�u�>�)����+��������ʦ�!�!�u�d�w�5�������� U��V��]���4�&�%�'���}�������]��y�����u�u�u�o�>�)����C����lǻ�����&��0���/����Y�ƿ�W9��P�����:�}��8�6�.�FϺ�����O��N�����u�&�:�3�3�/�W���Y����G��X	��*���!�'�d�1� �)�W���s�ƿ�T�������4�4�u�u�w�g��������l��C��D���:�;�:�e�l�}�����ƿ�	��^ �����u�u�u�!��2����������Z#����1�"�!�u�~�W�W��Y����R
��Q�����;�;�u�0� �8�W���Y����9F��N��1����4�;�!�>�}����Yۍ��^+��DN�����u�|�:�u�#�����&����\� N�����u�|�_�u�>�3�ϭ�=����[��N��U���!��4�9�)�M�������@[�X����r�r�|�_�w�$�ϟ�����Z�������,�}��8�6�.��������	��D�����6�#�6�:��}�������9F��^	��ʦ��1��4�9�}�W���Y����p��Y1��O���:�=�'�h��)����G���]ǻ��ʔ�6�8�=�<��}�Ͽ����X(��z��U���;�:�e�u�1�.��������V��EF�U���;�:�e�n�w�.����Y����P��_��U���u�u�6� ��<����C����G��DS����'�h�r�r�~�W�W�������@"��V8�����4�;�o�&�3�1��������AN��B�����:�;�:�e�w�`�_������V�d�����4�u�&�0�?�4�W���Y�����h�����0�!�'�>�"���������V�S�����'�h�r�r�l�}�����ƿ�r��Z8�����!�u�u�!��2����������Z#��ʱ�"�!�u�|�m�}�������A�=d�����4�u�&�4�6�<����Y�����h�����h�r�r�_�w�4����
����R/��N��U���o�&�1�9�0�>����������Y��E���h�}�!�0�$�c�G���s�ƿ�T������� �4�0�u�w�g��������\�^�����<�;�9�&��3�������F��D�����6�#�6�:��j��������\������k�e�|�_�w�4����
����|��T��U���o�&�1�9�0�>����������Y��E���h�}�!�0�$�c�G���s�ƿ�T�������9�1� ��;�g��������\�^�����<�;�9�&��)�!�������F��D�����6�o�u�e�l�W�W�������v��[������u�o�7�8�8���Y����V]ǑN�U���%�:�u�=�w��W���Y�����������1�!�0�u�2�3�W�������Z��C�����'�u�x�u��}��������G����ʱ�!�u�<�u�?�}�&ϼ����F��C�� ���>�0�u�u�#�4��ԜY����Z��RN�����3�&��!��1����Cӕ��]��^�����w�_�u�!�%�?��������UF��s��<���u�<�;�9�>�}����[����V��=d��Xǣ�:�>�0��9�������ƹK��_��*����&�!�3�;�8�Wύ�����]����U���<�,�"�'�y�$��������KF��c"��U���%�'�u�4�w�W�W���Y����V�N��H���4�&�y�u�w�}�W������\	��V ךU���u�4�%�0�;�}�W���*����V%��N��U���<�u�&�1�;�:����Y����R��R-��F���k��8�9��6����T�ƥ�F��S1�����u�u�u�&��(����Y���@��B ��U���u�x�u� �w�3��������\��XN����u�u�&�4�'�8�W���Gӕ��R��RG�U���x�:�!�7�8�8��ԶY����[	��h�����3�:�1�'�w��4���5����A��R �����:�>���2�����Y۴��l�N�����6�8�%�}�w�}�Wϵ�����@F������&�u�x�u�9�}��������W��N�����u�4�u�_�w�}�W���	����XF�N��Kʆ�8�9��>�w�}�W���Tӏ����h���ߊu�u�u�4�'�8����Y���F��Z��6���-�u�u�u�z�4�Wϭ�����ZǻN��U���4�%�0�u�w�}�J���
����_�N��U���x�<�u�7�8�8����Y����p	��{��U���u�h�u��2����Y���K�^ �����9�2�6�u�w�}�������F�N��U���0��y�u�w�}�W��Y���@��[�����u�u�&�:�1�4�W���Y�����R�����u�u�u�x�w�3�W���&����P9��T��]��1�"�!�u�~�}�W���
����U'��EN��U��u�&�:�3�3�/�W���Y���\��D�����6�#�6�:��}�������F�N��6�����'�,�w�c��������A��N��X��� �u�!�
�8�4�(�������}��V��Dʱ�"�!�u�|�w�}�Wϭ�:����R��N��H���&�:�3�4�6�}�W���T�ƣ�GF��S1�����#�6�:�}�`�9� ���Y��ƹF������;��0�&�j�}��������\��U��Xʺ�!�&�1�9�0�>�����Χ�F��T��U���;�:�e�_�]�}�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���l�C�����=�&�u�3�#�8�$������� �E�����u�:��8�;���������@F��X��U���x�u�4�0�"�1�[ϭ��Ƹ�R��_�����u�6� � �6�2�W���	����R��RN�����1�1�'�6�;�}�W��Y����[��V�����u�:�4�:�3�<�W�������R
�N��U���0�<�0�&�6�8�W�ԜY���K��_�����u�$�4�f�w�8����
Ӓ��GF��RN�����:�u�&�4�6�3����
����R0��^
��U���x�u� �!�5�}����Y����\��_��U���u�<�=�&��9�4������F��`�����e�u� �!�]�}�ZϮ�������ZN��U���4�%�0�_�w�p�W��Y���F�N��U���u�u�
�u�w��W���&���l9�N��U���
�u�u�
�w�}�(���Yӹ��l�C�����0�9�u�-�w�}�(���������KN��*���u�
�)�u��!�W����ư�l�K1��Uʩ�
�u�x�u�w�}�W���Y���F��h1��*���
�
�
�
���(���Y����l9��h1��*���
�
�
�
���(���T�ƿ�w��~ ��U���u�
��
��!�(���&�Ǝ�l9��h1��*���
�
�x�
���(���&����%��=N��X���u�u�u�u�w�}�Wρ�&����l9��h1��*���
�
�
�
�w�}�W���Y���F�1��*���
�
�_�u�z�.�3���/����z�N��U���u�u�u�u�w�}�W���Y�ư�l9��h1��*���
�
�)�u�z�W�W��
����A%��^ ��\���u�u�g�u�w�m�W���H�ư�T�KN��Uʩ�u�u�)�u�w�!�W�������ǻC�U���u�u�u�u�w�}�W���&����F�N��U���
�
�
�u�w�}�W���Yӹ��l9ǻC�����4�;�e�w�}�(���Y����l9��h1��*���u�u�u�
���(���&���F��h1��*���
�_�u�x�w�p�W��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���9lǻC�'���&�0�u�=�w�<�Ͽ�Ӑ��Z��Y��ʡ�u�#�<�u�6�:�W������@��RN�����u�x�u�<�9�1�W���ӄ��@��[�����=�u�-�1�:�4�W�������r%�:�����&�4�w�0�'�}��ԜY����[��^	�����:�u�=�!�%�<����ƭ�\��C��U���;�u�0�2�3�*�����ƥ�C��N�U���4�:�u�=�w�)��������	��C��U���!�'�_�u��:����
���C��R��&���9��>�-�]�}����s���Z ��^�����2�}�4�%�2�1�D�������F�N��U���:�;�h�d�u�)��ԜY���F��s��<���h�&�4�4�9�W�W���Y�ƿ�w��a�����i�u��!��1����s���F��SN��N���u�0�1�<�l�}����	����@��R	�����n�_�u�9��(��ԜY����V��d�����>�-�_�u�2�4�}���Y����Z��P1�����4�%�0�9�d�t����s���F�������h�e�w�!�2�W�W���Y�ƿ�d��V��E���h�r�r�_�w�}�W������F������<�}�|�i�w�m�L���Y����]��QUךU���;�u�3�_�w�3�W�������w
��X��N�ߊu�x��<�2�)�Ϸ�	����Z��[��ʡ�0�6�4�;�8�}�6���Yӕ��R��_��]���i�u�&�4�6�3�}���
����e��S-�����|�i�u�&�6�<����0��ƹ��T��6���;�e�u�h��)����G���l�D�����4�;�e�u�j�.��������V��EF��6���!�n�_�u�z�}����Y����}��V��Dʘ�� �<�&�]�}������ƹ ��'����!�u��8�6�.�FϹ�����VlǻN��X���:�
�u�$�6�n�}���Y�˺�\	��VN�������4�;��m�W���Tސ��\�������0�&��0� �����0���F�A�����&��4�<�0�2����
����Z��X��]���u�u�x�#�8�6�ϭ�=����]F��s��6���;��_�u�w�p����&�ƿ�w��x�����!��4�;��l�}���Y�˺�\	��VN��1����9�1�;�$���������R��~GךU���x�=�:�
�w�.��������F��D*�����<��4�;��l�}���Y�˺�\	��VN��1�����u�&�2�5����P���K��_��*���&�4�4�0�"�}��������zM��=N��U���=�:�
�u�$�9����0�ƿ�r��t���_�u�u�x�?�2�(���
����V��B�����'�=�<�}�|�t�W���Tސ��\��������u�&�6�"�����0���F�A�����&��6�8�"�}��������Z��_��U���x�#�:�>�6�.�6�������W)��������9�1� ��t�W���<���� �������"�'�{�$�6�n�Wǌ�5���F�P�����8�%�}�u�w�}�Wϵ�����]%��^ ��Kʜ�e�u�x�u�9�}�������� ��DךU���u�:�!�8�'�u�W���Y����R��R-��F���u�u�k��:�1�4������F�N��U���<�u�&�1�;�:����Y�����X�����u�u�u�k�$��������F�N��U���x�<�u�&�3�1��������AN��S�����|�u�u�u�w�.�4���.���F�S����0���'�.��[���Y���F��N�����2�6�u�u�w�}��������RF�N��Kʦ��0��!�{�}�W���Y���K�^ �����9�2�6�#�4�2�_������\F��=N��U���u�&�:�1�9�����Y����@*��S��6���&��y�u�w�}�ZϷ�Yӕ��l
��^ךU���u�u�&�4�6�3�W���Y�����V�����}�|�u�u�w�}�W������G��X	��*���!�'�d�u�8�3���s���F�D�����!�u�u�u�j�}��������]N��G�U���u�x�u� �w�)�(�������P��_����!�u�|�u�w�}�Wϭ�=����R
��~ ��U��&��!��;�9����Q���F�N��Uʦ�1�9�2�6�w�}�W���
����R0��^
�����k�&��!��1�����΅�O�C����&�1�9�2�4�}�W���Yӕ��R��R'��U���u�k�&���<�Ǘ�U���F�N��Xʼ�u�&�1�9�0�>�W���Y����@"��V9�� ���u�u�k�&� �����0���F�N��U����!�&�1�;�:����Y�����S
�����u�u�u�k�$���������J�N��U���x�<�u�&�3�1��������AN��S�����|�u�u�u�w�.�6�������GF�S����1��4�;��l�[���Y���F��CN�����2�6�#�6�8�u�W������l�N��Uʦ��6�8�;�w�}�W��Y����P��_��]���u�u�u�u�z�}��������T��A�����b�1�"�!�w�t�W���Y����@'��B�����u�u�k�&��>�����΅�O�N��U���:�!�&�1�;�:��������Q��X����_�u�u�u�w�.����/����|��
P����� ��9�1�"�u�^��Y���	����*���<�_�u�0�3�:�����Ƌ�]+��DUװ���x��<�u�$�)�ϸ�����P��B�����=�!�&�8�w�-�DϽ�����D	��_N��U���4�4�1�_�w�p��������RF��Y	��U��� �!�u�:�w�<�ύ�����_��N��[���=�&�<�u�$�3�W�ԜY����`6�������1�!�8�;�w�/����
Ӈ����RN�����9�2�6�u�w���������_��ETךU���6�&�}�4�'�8����P����V��=N��U���'�&�;�
�3�8�$������� �C�����u�u�&�6�"�(����E�Ƣ�GF��`�����>� ��6�~�W�W���Y����G��[�� ���h�&��6�:�<����ۍ��^+��DC�N���u�0�1�<�l�}����	����@��^ ��4���8�9�!�'�]�}�Z¨�����#��D����x�=�:�
�w���������]F��[��U���#�:�>�4��6�$������� ǻC�����
�u��}�#�8����I��ƹK��_��*�����u�d�]�}�Z�������P#��N��R���x�#�:�>�6�>�WǱ�����A��d��Xǣ�:�>�4�6�4�3��������R��\ ��8���|�u�x�#�8�6�Ͻ����l�C�����4�6�6� �w�-����Tސ��\�������;�9�6� �]�}�Z�������P#��������9�1� ������
���F�A�����6�6� � �6�8��������R��N��1���m�o�0�!�#�}����<����^�e:�����u�0�0�<�w�<�W�ԜY���X ��D��6���;�h�u�4�$�t�W������\	��V ��Hʳ�9�0�u�u�'�/�W���Y���F�t��U���u�u�h�u�6�-����J���F�N��U���u�u�x�u�9�}��������F�N��U���u�u�u�h�w�2����D����J�N��U���u�u�u�x�w�3�W���&����P9��T��]��1�"�!�u�~�}�W�������F�N��K��r�u�u�u�w�}�W���Y���F�N��Xʼ�u�&�1�9�0�>�W���YӅ��rT�N��U��r�r�u�u�w�}�W���Y���F�N��U���<�u�&�1�;�:����Y����qF�N��U���k�}�!�0�$�c�G���Y���F�N��U���x�<�u�&�3�1��������AN��
�����e�_�u�u�w��:���Y���X�I�U���u�u�u�u�w�}�W���Y���K��YN�����:�<�_�u�w�}�'���Y���F�������6�8�u�w�}�W���Y���F���U���
�:�<�
�2�)���Y����G	�d��U���6�;�u�u�w�}�J���
����^0��^
��¾� ��6�x�~�}�Z����ƿ�W9��P��U���u�6�6�;�w�}�W��Y����P��_��]���8�4�&�y�w�}�W��Y���@��[�����6�:�}�b�3�*����P���F��g�����u�u�k�:�2�q�W���Y���F�N��U���u�u�x�:�#�.��������V��EF�U���;�:�e�_�w�}�W�������R��
P����� � �4�0�l�}�W���Y���F�C�����!�
�:�<�]�W�W��-���� ��DN�����:�0�!�0�3�)�W���Ӓ��G��d�����>�1�8�<�{�*��������]ǻC����<�0� �u�2�;����Y����WF����U���&�u�3�!�2�����:������CN��ʠ�0�_�u�x�#�}��������R��^ ��U���u�<�!�'�4�<��ԶY���f��PN��1���%�3�'�!�2�8�����Ư�^��R ��U���!�4�u�u�6�}��������_	��=N��Xʰ�4�9�u�:�w�(����Ӫ��w��E�����!�u�;�u�1�8� ���
ӓ��Z
��Y�����4�<�<�,�w�p�W���Y����G�������'�:�!�:�w�5�W�������[��dךU���4�9��!�"��W��
����Q
��B�����r�r�_�u�z�����?����F�G������8�9��<�W�W�������F�C��U���<�2�0�2��<��������[��N��U���&�4�4� ��1�K�������T��A�����&�<�4��4�0�L���Y�����C����� ��9�i�w�.��������F��N��Xǰ�1�<�n�u�z�8�Ϯ�����)��G��3��_�u�0��#�(�1���Y����\�������;�9�6� �p�<��������GǻN��X���:�
�u��8�}��������9F�C�����
�u��&�#�<�W��s���K��X��ʴ�0�0�u�4�$�W�W���T����X9��T+�����7�0� �%�#�;�W���Tސ��\��-��U���%�0�9�_�w�}�Z�������P"��D(�����6�8�<�_�w�}�Z�������P7��s��:���6�}�|�u�w�����=������^�����{��:�u�%�1�}���Y�ƫ�]��TN�����u�u�u�u�<�8�������V�N�U���u�!�
�:�>�}�J���^���F��X�����}�u�u�u�w�<����Y����R
��N��U���u�u�u�x�>�}������ƹF�N��0���u�h�u��6�1�8�������F���U���9�4�_�u�w�}�W���Y���F��Z��6���u�u�u�u�z�}��������T��N��U���6�u�u�u�i�.�1�������^N��N��Xʼ�u�&�1�9�0�>�W���Y����bF�N��U���!��!�6��t�L���TӉ����h�����h�>�0�0��1�}����ƫ�]��C�����!� ��&�]�}�Z¨�����"��X�� ���!�4�4�4�>�W�W�������RF��R��#���r�r�u�x�!�2��������GF��[��U���#�:�>�4�4�3��������G��qךU���=�:�
�u�;�}��������F�A�����6�u�&�4�6�<���������X��U���&�4�4�4�>�����s�ƃ�G��s��#���1�u�;�<�.�*����?������d��Uʲ�;�'�6�8�'�u�W���YӍ��@��V��K��r�u�x�u�9�}��������	[�IךU���:�!�8�%��}�W�������GF������u�u�u�u�w�}�Z����Ʈ�\
��Yd��U���6�;�u�u�i�.��������F��N��X���;�u�:�9�6�W�W���Y����F�	N������>�u�u�w�}�W������G��X	�����u�u��u�w�`�W�������_��B�U���x�<�u�&�3�1����Y�����N��H����!��9�3�(�;���B���\��D�����6�o�u��$�)��Զs�ƿ�R��B��Hʦ�4�4� ��;�W�W�������Z��CN�U���!��9�1�"���Զ����g*��