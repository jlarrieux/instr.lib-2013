-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����J��X�����{�=�_�x��)���=����R��=C�:���<�4�u�'�=�>�Mύ�����K��X������u�x�u�6�8�W�������VǶd�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�}����I����\��^	��U���<�;�9��$�/����
ӥ��C	��C������9��2�#�}������ƴF��C�����;�!� �0�#�}��������] ��Z���߇x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�}��T�Ɯ�A��RT�����6�8�:�0�#�4��������RF��B ��ʡ�4�u�0�&�.�(��������IǶN��U���u�u�4�4�#�}�W��������������u�x�u�x�]�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���lǑ[�����<�0�n�u�"�8����W����_	��T1�C���9�n�u� �2�4��������P9��S@���ߠ0�!�!�u�.�>�����մ�Z�=���ߊu��&�!�w�}�W���Ʈ�\
��YUךU���%�0�9�u�w�g��������T��=N�����0�9�f�u�m�4�W���&����P]ǻ�����u�u�u�o�8�)��������F��@ ��U���_�u�&�4�'�8�W���CӉ����[��\���;�u�,�6�8�3����B����A��C�� �����:�u�.�>�����մ�ZǑN�����u�&�:�;��1�W���Y����T��_�����:�e�u�h�u�m�L���
����_F��X	�����u�u�o�7�8�8���Y����V]ǻ�����&��2�9��}�W������R�
N�����_�u�<�;�;�.�#�������V
������u�h�3�9�2�W�W�������@5��G�����u�u�:�9�6�}�Jϸ�����9F��C�����u�0�%�o�$�/���YӇ��A��C�����:�u�&�:�9���������������_�u�!�'�5�)�W���&����F��D����u�4�!�<�"�8��������GF����:����9�o�&�0�<�W���[���9l��P�����x��0�!�w�2����?���g���� ���u�:�&�:�w�5��������p
��R
��U���<�_�u�x��0��������\��Yd��!���9��o�u�'�2����*����V%��N�����0�<�u�u�w�W�W���Ӕ��Z��R
��]���%�0�9�|�#�8�}���Y�ƥ���D�����_�u�u�u�w�	����?��� ��D�U���u�0�&�_�w�}�W���-����V ��S������2�9��l�}�W�������U]ǻN�����3�_�u�;�w�/����Y����_��dךU����4�&�'��:����?Ӊ��AF��=�����9�f�u�:�6�3�W���Y����G	��R��U���;�0�_�u�8�3���YӖ��P��=�����9�f�|�<�]�}����s���Z ��^�����2�}�4�%�2�1�D�������F�N��U���&�!�!�0�]�}�W���Y����T��q��U��u�4�&�n�w�}�W���
����T
��Q*��U��3�9�0�_�w�}�W���
����G*��N��I���e�w�u�u�w�}�Wϭ�*����V*��N��Hʳ�9�0�_�u�w�}����Y���F�N�����9�6�u�:�6�3����
����@��[
��ʽ�;�9�1�%�8�8���� Ӓ��>��^ ��U���u�u�x�u�8�1�[ϼ�������NN��ʧ�9�!�1�6�8�6�������Q	����ʺ�!�:�u�u�w�}�W��Y����+��zG�U���u�u�&��0�1�1���Dӕ��T��q�U���u�u�&��0�1�1������@��P	��3��u�u�u�u�>�}��������w��O�����2�9��u�?�3�W���Y�����X��9���i�u�e�w�]�}�W���Y�ƿ�`��[����u�'�0�_�w�}�W�����ƹF�N��U���:�;��9�k�}��������M�d��U���u�u�&��:�1�;���E�ƪ�_��=N��U���u�;�u�3�]�}�W����ƥ�l�N��ʼ�n�u�0�1�'�2����:����V��=N�����;�u�h�&��(����B����@5��G��I���&�4�%�0�4�f�}���Y����9lǑ=d