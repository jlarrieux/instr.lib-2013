-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����A��s�����0�:�,�#�3�p�W�������y	��/�����;�x�u�'�0�3�ώ�����	F��~��C���_�x��!�m�o�W��� ����l�=C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�_�z�u�^��H�Ə�C��P��;���:�4�u�;�#�(����Y����\��^��X���9�u�<�=�$��������(��^��ʜ�&�'�8�;�$������ƅ�U	��V�����x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z�ԑTӶ��C	��N�����3�9�u�'�6�8�W���Y������X�����!�0�3�4�#�2��������G	��=C�U���u�u�u��>�}��������Z��E��U���d�g�u���<�ϫ��ƾ�R��E��U���;�0�&�x�w�}�W���Y�Ƹ���RN�����0�:�,�7�?�+�W���Ӈ��R��U�����!�u�=�3�w�8�������K�N��U���u��!��w�.� �������\F��RN�����0�:�,�4�3�8�ϩ��ƿ�R��Y8���߇x�u�u�u�w�}�������K�N��U���u�u�u�u�w�}��������W��D�����0�u�&�:�;�}�����ƻ�V��b�����4��1�0�$�p�W���Y���F��������0�%�<�#�/����������_N�����1�'�&��w�5����T���F�N�����1�0�1�1�%�.�>���
����@J��C�����u�!�<�u�2�/�������9K��C��U���u�u�u��#��Ϸ�Y����W����ʢ�&�'�4�u�%�0������ƴl�N��U���u�u��4��9�����ƥ�����ʴ�1�0�&�!�6�}����ӄ��@�������_�x�u�u�w�}�Wϰ��Ƽ�\��D��U���!�_�x�x�w�}�W���Y�Ƙ�VF��G�����0�4�u�'�:�.��������W��D'�����&�%�4�0�2�9����
���F�N��U���;�u��4��9����Ӓ��@"��V!��U���`�6�:�>�4�>���T���F�N��U���=�u�<�0�>�8���� Ӏ��^F��X�����1�'�&��w�3�W�������V��S
���߇x�u�u�u�w�}����
����r��R��ʡ�u��4��3�8����Y�����T�����{�x�_�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T����Z��E�����u�:�>�_�w�.�W���ݕ��l
��^��D��4�9�_�u�$�}��������Z��C
����u� �0�"�%�s��������P%��Q�����&�4�9�_�w�}�����Ɗ�R��R�����8�'�u�&�]�}����s���R4��R��U���7�:�0�;�]�}�W���	����XF��^ �����:�<�n�u�w�W�W���+����d��R/�����u�o�<�u�8�1���Y���F�D"�����1�1�'�&��}�W�������R��N�����4�0�0�1�3�/����Y����\	��V �U���&�0�1�1�%�.�>���Y����]��Y��Lʱ�"�!�u�|�w�p�"��H���FǻN��1�����9�1�m�4�W�������9F�������o�<�u�>�3���Y����G	�U��Xʆ�m�d�u�u�$�<����Y�ƥ���Y��D���:�;�:�e�l�p�W��W���FǻN��1����!�u�u�"�}��������W	��C��\���x�u�d�{�]�}�W�������bF��X�����0�}�b�1� �)�W���Y���`W��d��Uʦ�0�1�1�'�$��������]��Y��Lʱ�"�!�u�|�l�}�Zϋ�I����V��q������!��8�%�f�}�������G��<��U����4�!�0��)�:����ƥ�9F�=N�����9�&�0�:�.�g�5���JŹ��	[�X�����k�}�!�0�$�`�W��P��ƹl�D������!���;�9����Y�Ʈ�\
��YN�U���&�n�u�u�$�:����=����]0��^
�����o�7�:�0�9�g�W���
��ƹ��Y�����4�;�<�0�m�.����Q����\��XN�U��}�!�0�&�j�}�G���Y���`W��N��G���_�u�<�;�;�.���� ����z���*���<�
�0�!�%�n�W������]ǑN�����u��&�!�%�)�6�������C������u�h�3�9�2�}�}���������^�����&�u�u�;�>�3�������\F��T��]���0�&�h�u�g�t�W��Y����Vǻ�����&�0�1�1�%�.�W�������V�
�����e�o�u�:�?�/�W���^���F�;�[��u�&�2�4�w���������c��T�����;�1�l�1� �)�W���D�Σ�[��S�R��n�u�x� �g�l�}���������V
�����&�<� ��2�g��������
F��@ ��U���u�x�u�d�y�m�W�ԜY����R
��e��1����!�o�&�3�1��������AN��
�����e�o�u�:�?�/�W���^���9F��^	��ʦ�0�1�4�4�"����Cӕ��l
��^�����'�f�u�:�9�2�G���D�Σ�[��S�R��n�x�u�d�y�}�W�ԜY����R
��e��1����!�<�0�w�}��������E��X��@ʱ�"�!�u�|�m�}�������A��U��Xʆ�m�d�-�g�]�}��������X��T�����2�_�u�x��.��������[�������u�'�u�:�w�8��������\��EN��ʦ�u�=�!�!�2�/����ӂ��RǻC����=�u�0�:�.�4�W������R��^��ʾ�0�u�3�&�2�8� �������V��^��U���;�9�<�u�#�(�U�ԜY����Z��RN�����3�&�0�1�3�/����	����Z��[N��Uȡ� �w�_�u�#�/����Y����	��D*�����4�<��%��}����ӏ����RL�Uʴ�!�<� �0�<�8�W���
����z��[�����o�&�2�4�w�.�U�����ƹ��E�����0�%�:�u��)�>���	����Z��[N��Uȡ� �w�_�u�#�/����Y����	��D<�����4� ��%�f�}����ӏ����RL�U���u�u�u�x�!�2��������Gl�C�����&�2�;�_�5�:��ԜY����Z��^ �����&�4�4�;�6�4�W�������\F��^��3ʶ�;�7�u�9�4�9����Ӓ��G��Z�����u�x�u�!�2�*�����ƾ�F��PN�����!�u�=�u�2�2�Ͻ�����R�������2�3�<� �2�}�W��Y������CN��U���u�'�4�<�0�)�Ͻ�	����\ ��_�����0� �0�3�9�2����	����@��e��Ɔ�8�9��>�]�}����s���Z ��e�����=�;�u�u�w�.��������W6��R/��Hʳ�9�0�_�u�w�}�3���0����Z��G��I���4�&�n�u�w�8��������T9��P�����0�9�|�!�2�W�W���Y����R/��V��%����i�u��#��!������F�D*�����4�<��%��a�W�������R
��d��Uʰ�1�<�n�u�2�9��������FǻC�%���9�;�u�=�w�����Y����R
��XN������&�6�;�5�}����Ӆ��@��XN��ʸ�8�'�y�u�z�}��������G��E�����1�9�,�!�w�5�W�������\�������u�<�<�2�1�4����Y����A	��D��'���!��8�9��6�}�������F�^��'���!�u�=�;�w�}�Wϭ�����c��R��]���0�&�h�u�g�t�}���Y����UF��D��*���0��8�9��6�W������F��s��<���%�u�h�&�6�<����Y����R/��d��Uʰ�1�<�n�u�2�9��������9F�-�����!�0��<�2�����
ӥ��]��=N�����&�}��&�#�����:���F��P��U���<�}��&�#�}����Y�����^�����&�u�h�}�#�8���Y���l�N�����0��<�0�3�/����	��� ��D�U���0�&�3�'�$�3�(���۵��C
��[�����_�u�u�u��.��������A��g��U��&�0�0��>�8����
��ƹF������0��<�0�3�/����	�Ƹ�VǻN��U����<�0�1�%�.�W��Q����A�	N��R��u�u�u�0�$�;��������_��^��\ʡ�0�u�u�u�w�}��������A��R�����!��1�0�$�v�F�ԜY���V��^�U���0�1�<�n�w�8�Ϯ�����l�=N��Xʖ�0�!�u�=�w�8�ϟ�����%��Y�����'�6�&�}��.�Í�����_�N�����u�u�<�}��.������ƹF������1�0�&�i�w�2����Y���A�=N��U���<�u�<�<�0�8��������p
�������u�u�<�}��9��������A�������u�u�u�<����������A��~ �����u�u�u�u�w�}��������V��S��'����1�0�&�9�W�W���Y�Ʃ�@ǻN��U���u��4��3�8���Y����W'��E��8���&�;�n�u�w�}�Wϻ�ӏ��9F�N�����3�_�u�u�9�}��ԜY����C��R�����u�&�0�1�3�/��������VF������1�0�&�x�f�W�W���T�Ɯ�C��Y������4��1�2�.�����ƿ���D��3���4�u�0�%�6�8�W���
�Ƹ��������_�u�x�:�?�/��������\��Y	�����u�:�!�0�:�0��������P��RN�����;�u�4�9�%�s�}�������@N��R��Y���%�0�9�|�w�?����Y����UN��R��\ʡ�0�_�u�u�w���������c��R��]���0�&�h�u�g�t�}���Y����UF��D��*���0��8�9��6�W������F��e��4���0�&�<�0�k�}�%���8����@��N�����<�n�u�0�3�-����
���Fǻ������!��u�j�.��������V��EF�����;�<�0�n�w�W�W��:����VF��RN�����_�u�x��;�2�W���Y����PF��SN��ʦ�:�9�u�0�>�-��������@F��XN������_�u�%�>��������p
��=N�����_�u�u�3�%�.��������R��R-��\ʡ�0�_�u�u�w�;��������_��^��\ʡ�0�u�u�u�w�}�Wϭ�������^ �����&�'�!��3�8����E�ƿ�V��N*�����_�u�u�u�9�}��ԜY���@4��S*�����u�h�&�0�8�$��������AN��R�����&��%�|�l�}�W���
����w��x�����u�h�&�0�3�<����B����������;�u�'�6�$�f�W�ԜY����Z��^ �����1�!�u� �'�)��������Z��PN�����:�8�0�u�2�*�����ơ�^	��=N��Xʴ�1�!�0���W�W�������R4��R�&���9��>�_�w�8��ԜY�ƥ���D��U���;�u�u�u�$�8��������Z��R��]���0�&�h�u�g�t�}���Y����UF��D��*���0��8�9��6�W������F��e��1����!�<�0�w�`��������|��^��N���u�0�1�<�l�}����	����@��N�����x��&�2�w�5�W���	����F��V�� ���i�u�<�;�3�.��������G6��R_��@ʱ�"�!�u�m�~�W�W�������bF������&�0�1�4�6�(�'���H����W	��C��\��u�&�0�1�3�/�������@4��S/������;�&�;�l�}�W����ƞ�]�