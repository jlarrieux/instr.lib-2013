-- � 2012 National Instruments Corporation.
encrypted

�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�W�ZϘ�����B%��Q"�����#�1�x�u�"�5�����Ǝ�X��C�����;�9��:�2�)�W�������4ǶN����g�u�4� �%�}�G��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�u�6�u�g�l�4�������(��^��ʜ�&�'�8�;�$���������9K�v��'���!�u�0�0�!�9�Z�������R
��Y�� ���!�u�;�0�9�1�>�������\ǶC�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�_�x�z�}����
����[��T�����!�!�>�&�>�}��������P��CN�����<�;�9�y�6�9��������K������ �9�&�2�6�.��������\ ��_��4���_�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T���K�C�X���x�x�x�x�z�p�Z��T����Z��E�����_�u�&�u�2�8��������lW��@���ߊu�&�u�0�2�3����������d�����,���0��<����
����V��^��Uʾ� ��6�u�w�}�W���ӏ��V��T��D���n�%�'�}�w�����:���F�N��U���
�:�<�n�w�����:����F�N��U���
�:�<�n�w�.�$������F�N��U���9�4�n�_�w��������F������9�2�6�_�w�����Y���F������9�2�6�_�w��������F������9�2�6�#�4�2�_������\F��dךU���:�3�1�'�w�}�Mϱ�ӕ��l
��^�����'�d�1�"�#�}�^�ԜY����V ��v�����u� �u�!��2����������Z#����1�"�!�u�~�W�W�������G�N��U���u�!�
�:�>���������W	��C��\�ߊu�&�:�1�9�����CӉ����h�����0�!�'�>�"����Y����G	�N����u�$�:�3�8�9��Զs����Z��C��U���u�3���2�����Y��ƓF�=�����=�'�u�<�;�?�W���Ӊ��G��RN��U���u��3�9�2�q����[������XNךU���0�&�'�u�?�$����Ӂ����P�����!�0�u�;�w�<����������B��Uʦ�2�4�u��2��������\��C
�����u�h�r�r�]�}����ӕ��V ��e��U���u�o�&�1�;�:���Y���9F��^	��ʦ�:�3�<��0�}�W���Y����_	��T1�����}�b�1�"�#�}�^��Yۉ��V��	I�\�ߊu�<�;�9�$���������F�N�����0�}�u�:�9�2�G���D�Σ�[��
P��R��u�&�2�4�w�.�������F�T�����:�<�
�0�#�/����4����F��@ ��U���o�u�:�=�%�`�P���B����Z��[N��6����!��9�w�}�W���&����P9��T��]��1�"�!�u�~�g�WǱ�����A��UךU���;�9�&��2�
�6��� ����	F��S1�����#�6�:�}��0����Hӂ��]��G��H���!�0�&�k�g�t�}���������X�����u�u�u�o�$�9�������V�=d�����<� �0�>�2�}�W�������F��C�� ���>�0�u�3�$�2��������F�N�����u�&�w�'�2�f�WϿ�����G��R������0���0�}�W���Cӕ��]��^�����w�_�u�!�%�?��������UF��X�����2�u�u�u�w�4��������A��d�����<� �0�>�2�}�ϭ�:����\��R��U��&�2�4�u�$�����B����G��U��U���%�:�u�&�2�5����Y���\��^	��ʼ�u�!� �w�]�}��������X�������0��!��;�}�W�������������u�4�!�<�"�8����Y����@%��Q9������9�o�&�0�<�W���[����]ǻ�����!�u�0�%�8�}��������JF�N��U���;�9�<�u�#�(�U�ԶYӇ��A��C�����4�:�!�u�#�4��ԜY����Z��RN�����;� �u�3�$���������\��^	��ʼ�u�b�n�u�6�)����Ӌ��l ��X�����&�:�3�4�6�>�W���������Y����2�;�_�u�z������ƭ�_F��G��U���%�:�0�!�6�<��������]��E��U���<�u�;�!�2��}���Tӂ��T��N�����w�:�u�=�$�}�����Ƹ���^
�����;�"�!�u�?�}����Y���F��[��ʼ�u�=�u��!�s�W���
Ӈ��@F��(��ʺ�0�4�9�!�w�5�W�������bl�C�����'�u�;�u�"�)���� �Ƹ�VF��V
��ʺ�u�=�u�:�1�4����
ӄ��F��T�����0�<�!�'�;�����C����A	��D�����0�9�|�u�5�:����Yӏ��A��Y	������8�9��<�}����Y�����R�����2�i�u��2����Y�����R��'���i�u��0� �f�W���Yӕ��V ��Y<��U��&�:�3�<�l�}�Wϻ�ӏ��9F��Y
�����&�u�0�<�#�/����	����9l�C�����6�1�u�:�9�.� ���Ӆ��U ��^��U���'�u�;�}�z�t�W���Y����RF��^��U���u�0�<�!�%�)�W���	Ӓ��P��QN�������"�r�2�2�Wǭ�.����U�=d��X�����u�=�$�-����
Ӆ��_��V�����u�;�!�0��0����ӂ��R����U���<�2�u�x�w�2�$������� ��^�����9�u�3�&��0����Ӓ����V��ʦ�8�u�d�&�w�p�W�������R��E�����u�<�<�-�w�5�ϗ������������u�:�!�0�#�2�ϰ����F��X�����:�%�!�;�w�5�W���
�ƨ�U ��R ��U���"�0�u�=�w�1��������@Hǻ/������ �!�'�]�}����
�Ο�^��t���ߊu�0�<�_�w�}�Ϭ�
����V��=�����9�f�|�!�2�W�W���Y����@5��G�����_�u�u�u�w�4�W�������W4��
I�U���;�u�u�u�w�}��������]��R��]���0�&�k�e�~�W�W���Y���@��d����u�:�=�'�j�z�P��Y���F������3�}�|�i�w�l�L���Y�����^��6�����2�r�p�)��ԜY���F�^�����3�:�;�0�j�l�UϪ����F�N��Uʦ��0�� �#�/�K�������@[�I����u�u�u�u�w�.���������R=������8�4�&�e�9� ���Y���A��d��U���u�u�0�&�]�}�W���Y���@��R�� ���'�i�u�&�8�;�������]ǻN��U���u�;�u�3�]�}�W���Y����Z ��=N��U���;�u�3�_�w�}�������V��G������1�0�&�8�3���s�ƿ�p	��v
��U��&�1�9�2�4�+����Q����V ��B ����_�u�x��>�}����������^�� ���"�<�0�0�6�1�ϸ�Ӄ��[F����U���&�u�=�6�w�}�Z�������[����U���u�,�9�u�8�}��������Z��YךU���%�!�0�o�w�-����
۵��C
��[��\���7�2�;�u�w�4�W�������W��d�����>�-�u�=�9�}�W���
����U1��[��Hʦ�:�3�0�0�l�}�W���������N��U���8�4�&�d�;�2�}���Y���@��R��4���,�6�}�|�k�}��������zO��Y
��6�����2�4�3�3�ϭ�:����V"��d��U���0�1�9�:�l�}�W����ƿ�\��R<��H��u�=�;�u�w�}�Wϭ�:����R��T��Hʦ�:�3�<��0�W�W���Y����Z ��N�����<�n�u�0�3�-����
ө��C��R����&�:�3�4�6�a�W�������G��[UךU���:�3�0�'�6�}�Jϭ�:����V'��V���ߊu�&�:�1�9�����E�ƿ�d��^����1���_